module clock(output clock_signal);

(* LOC="Y19" *) IB clock_pin(clock_signal);

endmodule
