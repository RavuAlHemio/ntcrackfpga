module state_giver(
    input clk,
    input [4:0] password_len,
    input [159:0] password_chars,
    input [(128*128-1):0] hashes,
    input [127:0] current_hash,
    output reg [7:0] state_byte);

reg [11:0] byte_index;

initial begin
    byte_index <= 0;
end

always @ (posedge clk) begin
    case (byte_index)
        /* header */
        0: state_byte <= 8'h0A;
        1: state_byte <= 8'h55;
        2: state_byte <= 8'hFA;
        3: state_byte <= 8'hCE;

        // password length
        4: state_byte <= password_len;

        // password characters
        5: state_byte <= password_chars[159:152];
        6: state_byte <= password_chars[151:144];
        7: state_byte <= password_chars[143:136];
        8: state_byte <= password_chars[135:128];
        9: state_byte <= password_chars[127:120];
        10: state_byte <= password_chars[119:112];
        11: state_byte <= password_chars[111:104];
        12: state_byte <= password_chars[103:96];
        13: state_byte <= password_chars[95:88];
        14: state_byte <= password_chars[87:80];
        15: state_byte <= password_chars[79:72];
        16: state_byte <= password_chars[71:64];
        17: state_byte <= password_chars[63:56];
        18: state_byte <= password_chars[55:48];
        19: state_byte <= password_chars[47:40];
        20: state_byte <= password_chars[39:32];
        21: state_byte <= password_chars[31:24];
        22: state_byte <= password_chars[23:16];
        23: state_byte <= password_chars[15:8];
        24: state_byte <= password_chars[7:0];

        // stored hashes
        // Python:
        // for n in range(2048):
        //     print(f"        {n+25}: state_byte <= hashes[{128*128-(8*n+1)}:{128*128-(8*n+8)}];")
        25: state_byte <= hashes[16383:16376];
        26: state_byte <= hashes[16375:16368];
        27: state_byte <= hashes[16367:16360];
        28: state_byte <= hashes[16359:16352];
        29: state_byte <= hashes[16351:16344];
        30: state_byte <= hashes[16343:16336];
        31: state_byte <= hashes[16335:16328];
        32: state_byte <= hashes[16327:16320];
        33: state_byte <= hashes[16319:16312];
        34: state_byte <= hashes[16311:16304];
        35: state_byte <= hashes[16303:16296];
        36: state_byte <= hashes[16295:16288];
        37: state_byte <= hashes[16287:16280];
        38: state_byte <= hashes[16279:16272];
        39: state_byte <= hashes[16271:16264];
        40: state_byte <= hashes[16263:16256];
        41: state_byte <= hashes[16255:16248];
        42: state_byte <= hashes[16247:16240];
        43: state_byte <= hashes[16239:16232];
        44: state_byte <= hashes[16231:16224];
        45: state_byte <= hashes[16223:16216];
        46: state_byte <= hashes[16215:16208];
        47: state_byte <= hashes[16207:16200];
        48: state_byte <= hashes[16199:16192];
        49: state_byte <= hashes[16191:16184];
        50: state_byte <= hashes[16183:16176];
        51: state_byte <= hashes[16175:16168];
        52: state_byte <= hashes[16167:16160];
        53: state_byte <= hashes[16159:16152];
        54: state_byte <= hashes[16151:16144];
        55: state_byte <= hashes[16143:16136];
        56: state_byte <= hashes[16135:16128];
        57: state_byte <= hashes[16127:16120];
        58: state_byte <= hashes[16119:16112];
        59: state_byte <= hashes[16111:16104];
        60: state_byte <= hashes[16103:16096];
        61: state_byte <= hashes[16095:16088];
        62: state_byte <= hashes[16087:16080];
        63: state_byte <= hashes[16079:16072];
        64: state_byte <= hashes[16071:16064];
        65: state_byte <= hashes[16063:16056];
        66: state_byte <= hashes[16055:16048];
        67: state_byte <= hashes[16047:16040];
        68: state_byte <= hashes[16039:16032];
        69: state_byte <= hashes[16031:16024];
        70: state_byte <= hashes[16023:16016];
        71: state_byte <= hashes[16015:16008];
        72: state_byte <= hashes[16007:16000];
        73: state_byte <= hashes[15999:15992];
        74: state_byte <= hashes[15991:15984];
        75: state_byte <= hashes[15983:15976];
        76: state_byte <= hashes[15975:15968];
        77: state_byte <= hashes[15967:15960];
        78: state_byte <= hashes[15959:15952];
        79: state_byte <= hashes[15951:15944];
        80: state_byte <= hashes[15943:15936];
        81: state_byte <= hashes[15935:15928];
        82: state_byte <= hashes[15927:15920];
        83: state_byte <= hashes[15919:15912];
        84: state_byte <= hashes[15911:15904];
        85: state_byte <= hashes[15903:15896];
        86: state_byte <= hashes[15895:15888];
        87: state_byte <= hashes[15887:15880];
        88: state_byte <= hashes[15879:15872];
        89: state_byte <= hashes[15871:15864];
        90: state_byte <= hashes[15863:15856];
        91: state_byte <= hashes[15855:15848];
        92: state_byte <= hashes[15847:15840];
        93: state_byte <= hashes[15839:15832];
        94: state_byte <= hashes[15831:15824];
        95: state_byte <= hashes[15823:15816];
        96: state_byte <= hashes[15815:15808];
        97: state_byte <= hashes[15807:15800];
        98: state_byte <= hashes[15799:15792];
        99: state_byte <= hashes[15791:15784];
        100: state_byte <= hashes[15783:15776];
        101: state_byte <= hashes[15775:15768];
        102: state_byte <= hashes[15767:15760];
        103: state_byte <= hashes[15759:15752];
        104: state_byte <= hashes[15751:15744];
        105: state_byte <= hashes[15743:15736];
        106: state_byte <= hashes[15735:15728];
        107: state_byte <= hashes[15727:15720];
        108: state_byte <= hashes[15719:15712];
        109: state_byte <= hashes[15711:15704];
        110: state_byte <= hashes[15703:15696];
        111: state_byte <= hashes[15695:15688];
        112: state_byte <= hashes[15687:15680];
        113: state_byte <= hashes[15679:15672];
        114: state_byte <= hashes[15671:15664];
        115: state_byte <= hashes[15663:15656];
        116: state_byte <= hashes[15655:15648];
        117: state_byte <= hashes[15647:15640];
        118: state_byte <= hashes[15639:15632];
        119: state_byte <= hashes[15631:15624];
        120: state_byte <= hashes[15623:15616];
        121: state_byte <= hashes[15615:15608];
        122: state_byte <= hashes[15607:15600];
        123: state_byte <= hashes[15599:15592];
        124: state_byte <= hashes[15591:15584];
        125: state_byte <= hashes[15583:15576];
        126: state_byte <= hashes[15575:15568];
        127: state_byte <= hashes[15567:15560];
        128: state_byte <= hashes[15559:15552];
        129: state_byte <= hashes[15551:15544];
        130: state_byte <= hashes[15543:15536];
        131: state_byte <= hashes[15535:15528];
        132: state_byte <= hashes[15527:15520];
        133: state_byte <= hashes[15519:15512];
        134: state_byte <= hashes[15511:15504];
        135: state_byte <= hashes[15503:15496];
        136: state_byte <= hashes[15495:15488];
        137: state_byte <= hashes[15487:15480];
        138: state_byte <= hashes[15479:15472];
        139: state_byte <= hashes[15471:15464];
        140: state_byte <= hashes[15463:15456];
        141: state_byte <= hashes[15455:15448];
        142: state_byte <= hashes[15447:15440];
        143: state_byte <= hashes[15439:15432];
        144: state_byte <= hashes[15431:15424];
        145: state_byte <= hashes[15423:15416];
        146: state_byte <= hashes[15415:15408];
        147: state_byte <= hashes[15407:15400];
        148: state_byte <= hashes[15399:15392];
        149: state_byte <= hashes[15391:15384];
        150: state_byte <= hashes[15383:15376];
        151: state_byte <= hashes[15375:15368];
        152: state_byte <= hashes[15367:15360];
        153: state_byte <= hashes[15359:15352];
        154: state_byte <= hashes[15351:15344];
        155: state_byte <= hashes[15343:15336];
        156: state_byte <= hashes[15335:15328];
        157: state_byte <= hashes[15327:15320];
        158: state_byte <= hashes[15319:15312];
        159: state_byte <= hashes[15311:15304];
        160: state_byte <= hashes[15303:15296];
        161: state_byte <= hashes[15295:15288];
        162: state_byte <= hashes[15287:15280];
        163: state_byte <= hashes[15279:15272];
        164: state_byte <= hashes[15271:15264];
        165: state_byte <= hashes[15263:15256];
        166: state_byte <= hashes[15255:15248];
        167: state_byte <= hashes[15247:15240];
        168: state_byte <= hashes[15239:15232];
        169: state_byte <= hashes[15231:15224];
        170: state_byte <= hashes[15223:15216];
        171: state_byte <= hashes[15215:15208];
        172: state_byte <= hashes[15207:15200];
        173: state_byte <= hashes[15199:15192];
        174: state_byte <= hashes[15191:15184];
        175: state_byte <= hashes[15183:15176];
        176: state_byte <= hashes[15175:15168];
        177: state_byte <= hashes[15167:15160];
        178: state_byte <= hashes[15159:15152];
        179: state_byte <= hashes[15151:15144];
        180: state_byte <= hashes[15143:15136];
        181: state_byte <= hashes[15135:15128];
        182: state_byte <= hashes[15127:15120];
        183: state_byte <= hashes[15119:15112];
        184: state_byte <= hashes[15111:15104];
        185: state_byte <= hashes[15103:15096];
        186: state_byte <= hashes[15095:15088];
        187: state_byte <= hashes[15087:15080];
        188: state_byte <= hashes[15079:15072];
        189: state_byte <= hashes[15071:15064];
        190: state_byte <= hashes[15063:15056];
        191: state_byte <= hashes[15055:15048];
        192: state_byte <= hashes[15047:15040];
        193: state_byte <= hashes[15039:15032];
        194: state_byte <= hashes[15031:15024];
        195: state_byte <= hashes[15023:15016];
        196: state_byte <= hashes[15015:15008];
        197: state_byte <= hashes[15007:15000];
        198: state_byte <= hashes[14999:14992];
        199: state_byte <= hashes[14991:14984];
        200: state_byte <= hashes[14983:14976];
        201: state_byte <= hashes[14975:14968];
        202: state_byte <= hashes[14967:14960];
        203: state_byte <= hashes[14959:14952];
        204: state_byte <= hashes[14951:14944];
        205: state_byte <= hashes[14943:14936];
        206: state_byte <= hashes[14935:14928];
        207: state_byte <= hashes[14927:14920];
        208: state_byte <= hashes[14919:14912];
        209: state_byte <= hashes[14911:14904];
        210: state_byte <= hashes[14903:14896];
        211: state_byte <= hashes[14895:14888];
        212: state_byte <= hashes[14887:14880];
        213: state_byte <= hashes[14879:14872];
        214: state_byte <= hashes[14871:14864];
        215: state_byte <= hashes[14863:14856];
        216: state_byte <= hashes[14855:14848];
        217: state_byte <= hashes[14847:14840];
        218: state_byte <= hashes[14839:14832];
        219: state_byte <= hashes[14831:14824];
        220: state_byte <= hashes[14823:14816];
        221: state_byte <= hashes[14815:14808];
        222: state_byte <= hashes[14807:14800];
        223: state_byte <= hashes[14799:14792];
        224: state_byte <= hashes[14791:14784];
        225: state_byte <= hashes[14783:14776];
        226: state_byte <= hashes[14775:14768];
        227: state_byte <= hashes[14767:14760];
        228: state_byte <= hashes[14759:14752];
        229: state_byte <= hashes[14751:14744];
        230: state_byte <= hashes[14743:14736];
        231: state_byte <= hashes[14735:14728];
        232: state_byte <= hashes[14727:14720];
        233: state_byte <= hashes[14719:14712];
        234: state_byte <= hashes[14711:14704];
        235: state_byte <= hashes[14703:14696];
        236: state_byte <= hashes[14695:14688];
        237: state_byte <= hashes[14687:14680];
        238: state_byte <= hashes[14679:14672];
        239: state_byte <= hashes[14671:14664];
        240: state_byte <= hashes[14663:14656];
        241: state_byte <= hashes[14655:14648];
        242: state_byte <= hashes[14647:14640];
        243: state_byte <= hashes[14639:14632];
        244: state_byte <= hashes[14631:14624];
        245: state_byte <= hashes[14623:14616];
        246: state_byte <= hashes[14615:14608];
        247: state_byte <= hashes[14607:14600];
        248: state_byte <= hashes[14599:14592];
        249: state_byte <= hashes[14591:14584];
        250: state_byte <= hashes[14583:14576];
        251: state_byte <= hashes[14575:14568];
        252: state_byte <= hashes[14567:14560];
        253: state_byte <= hashes[14559:14552];
        254: state_byte <= hashes[14551:14544];
        255: state_byte <= hashes[14543:14536];
        256: state_byte <= hashes[14535:14528];
        257: state_byte <= hashes[14527:14520];
        258: state_byte <= hashes[14519:14512];
        259: state_byte <= hashes[14511:14504];
        260: state_byte <= hashes[14503:14496];
        261: state_byte <= hashes[14495:14488];
        262: state_byte <= hashes[14487:14480];
        263: state_byte <= hashes[14479:14472];
        264: state_byte <= hashes[14471:14464];
        265: state_byte <= hashes[14463:14456];
        266: state_byte <= hashes[14455:14448];
        267: state_byte <= hashes[14447:14440];
        268: state_byte <= hashes[14439:14432];
        269: state_byte <= hashes[14431:14424];
        270: state_byte <= hashes[14423:14416];
        271: state_byte <= hashes[14415:14408];
        272: state_byte <= hashes[14407:14400];
        273: state_byte <= hashes[14399:14392];
        274: state_byte <= hashes[14391:14384];
        275: state_byte <= hashes[14383:14376];
        276: state_byte <= hashes[14375:14368];
        277: state_byte <= hashes[14367:14360];
        278: state_byte <= hashes[14359:14352];
        279: state_byte <= hashes[14351:14344];
        280: state_byte <= hashes[14343:14336];
        281: state_byte <= hashes[14335:14328];
        282: state_byte <= hashes[14327:14320];
        283: state_byte <= hashes[14319:14312];
        284: state_byte <= hashes[14311:14304];
        285: state_byte <= hashes[14303:14296];
        286: state_byte <= hashes[14295:14288];
        287: state_byte <= hashes[14287:14280];
        288: state_byte <= hashes[14279:14272];
        289: state_byte <= hashes[14271:14264];
        290: state_byte <= hashes[14263:14256];
        291: state_byte <= hashes[14255:14248];
        292: state_byte <= hashes[14247:14240];
        293: state_byte <= hashes[14239:14232];
        294: state_byte <= hashes[14231:14224];
        295: state_byte <= hashes[14223:14216];
        296: state_byte <= hashes[14215:14208];
        297: state_byte <= hashes[14207:14200];
        298: state_byte <= hashes[14199:14192];
        299: state_byte <= hashes[14191:14184];
        300: state_byte <= hashes[14183:14176];
        301: state_byte <= hashes[14175:14168];
        302: state_byte <= hashes[14167:14160];
        303: state_byte <= hashes[14159:14152];
        304: state_byte <= hashes[14151:14144];
        305: state_byte <= hashes[14143:14136];
        306: state_byte <= hashes[14135:14128];
        307: state_byte <= hashes[14127:14120];
        308: state_byte <= hashes[14119:14112];
        309: state_byte <= hashes[14111:14104];
        310: state_byte <= hashes[14103:14096];
        311: state_byte <= hashes[14095:14088];
        312: state_byte <= hashes[14087:14080];
        313: state_byte <= hashes[14079:14072];
        314: state_byte <= hashes[14071:14064];
        315: state_byte <= hashes[14063:14056];
        316: state_byte <= hashes[14055:14048];
        317: state_byte <= hashes[14047:14040];
        318: state_byte <= hashes[14039:14032];
        319: state_byte <= hashes[14031:14024];
        320: state_byte <= hashes[14023:14016];
        321: state_byte <= hashes[14015:14008];
        322: state_byte <= hashes[14007:14000];
        323: state_byte <= hashes[13999:13992];
        324: state_byte <= hashes[13991:13984];
        325: state_byte <= hashes[13983:13976];
        326: state_byte <= hashes[13975:13968];
        327: state_byte <= hashes[13967:13960];
        328: state_byte <= hashes[13959:13952];
        329: state_byte <= hashes[13951:13944];
        330: state_byte <= hashes[13943:13936];
        331: state_byte <= hashes[13935:13928];
        332: state_byte <= hashes[13927:13920];
        333: state_byte <= hashes[13919:13912];
        334: state_byte <= hashes[13911:13904];
        335: state_byte <= hashes[13903:13896];
        336: state_byte <= hashes[13895:13888];
        337: state_byte <= hashes[13887:13880];
        338: state_byte <= hashes[13879:13872];
        339: state_byte <= hashes[13871:13864];
        340: state_byte <= hashes[13863:13856];
        341: state_byte <= hashes[13855:13848];
        342: state_byte <= hashes[13847:13840];
        343: state_byte <= hashes[13839:13832];
        344: state_byte <= hashes[13831:13824];
        345: state_byte <= hashes[13823:13816];
        346: state_byte <= hashes[13815:13808];
        347: state_byte <= hashes[13807:13800];
        348: state_byte <= hashes[13799:13792];
        349: state_byte <= hashes[13791:13784];
        350: state_byte <= hashes[13783:13776];
        351: state_byte <= hashes[13775:13768];
        352: state_byte <= hashes[13767:13760];
        353: state_byte <= hashes[13759:13752];
        354: state_byte <= hashes[13751:13744];
        355: state_byte <= hashes[13743:13736];
        356: state_byte <= hashes[13735:13728];
        357: state_byte <= hashes[13727:13720];
        358: state_byte <= hashes[13719:13712];
        359: state_byte <= hashes[13711:13704];
        360: state_byte <= hashes[13703:13696];
        361: state_byte <= hashes[13695:13688];
        362: state_byte <= hashes[13687:13680];
        363: state_byte <= hashes[13679:13672];
        364: state_byte <= hashes[13671:13664];
        365: state_byte <= hashes[13663:13656];
        366: state_byte <= hashes[13655:13648];
        367: state_byte <= hashes[13647:13640];
        368: state_byte <= hashes[13639:13632];
        369: state_byte <= hashes[13631:13624];
        370: state_byte <= hashes[13623:13616];
        371: state_byte <= hashes[13615:13608];
        372: state_byte <= hashes[13607:13600];
        373: state_byte <= hashes[13599:13592];
        374: state_byte <= hashes[13591:13584];
        375: state_byte <= hashes[13583:13576];
        376: state_byte <= hashes[13575:13568];
        377: state_byte <= hashes[13567:13560];
        378: state_byte <= hashes[13559:13552];
        379: state_byte <= hashes[13551:13544];
        380: state_byte <= hashes[13543:13536];
        381: state_byte <= hashes[13535:13528];
        382: state_byte <= hashes[13527:13520];
        383: state_byte <= hashes[13519:13512];
        384: state_byte <= hashes[13511:13504];
        385: state_byte <= hashes[13503:13496];
        386: state_byte <= hashes[13495:13488];
        387: state_byte <= hashes[13487:13480];
        388: state_byte <= hashes[13479:13472];
        389: state_byte <= hashes[13471:13464];
        390: state_byte <= hashes[13463:13456];
        391: state_byte <= hashes[13455:13448];
        392: state_byte <= hashes[13447:13440];
        393: state_byte <= hashes[13439:13432];
        394: state_byte <= hashes[13431:13424];
        395: state_byte <= hashes[13423:13416];
        396: state_byte <= hashes[13415:13408];
        397: state_byte <= hashes[13407:13400];
        398: state_byte <= hashes[13399:13392];
        399: state_byte <= hashes[13391:13384];
        400: state_byte <= hashes[13383:13376];
        401: state_byte <= hashes[13375:13368];
        402: state_byte <= hashes[13367:13360];
        403: state_byte <= hashes[13359:13352];
        404: state_byte <= hashes[13351:13344];
        405: state_byte <= hashes[13343:13336];
        406: state_byte <= hashes[13335:13328];
        407: state_byte <= hashes[13327:13320];
        408: state_byte <= hashes[13319:13312];
        409: state_byte <= hashes[13311:13304];
        410: state_byte <= hashes[13303:13296];
        411: state_byte <= hashes[13295:13288];
        412: state_byte <= hashes[13287:13280];
        413: state_byte <= hashes[13279:13272];
        414: state_byte <= hashes[13271:13264];
        415: state_byte <= hashes[13263:13256];
        416: state_byte <= hashes[13255:13248];
        417: state_byte <= hashes[13247:13240];
        418: state_byte <= hashes[13239:13232];
        419: state_byte <= hashes[13231:13224];
        420: state_byte <= hashes[13223:13216];
        421: state_byte <= hashes[13215:13208];
        422: state_byte <= hashes[13207:13200];
        423: state_byte <= hashes[13199:13192];
        424: state_byte <= hashes[13191:13184];
        425: state_byte <= hashes[13183:13176];
        426: state_byte <= hashes[13175:13168];
        427: state_byte <= hashes[13167:13160];
        428: state_byte <= hashes[13159:13152];
        429: state_byte <= hashes[13151:13144];
        430: state_byte <= hashes[13143:13136];
        431: state_byte <= hashes[13135:13128];
        432: state_byte <= hashes[13127:13120];
        433: state_byte <= hashes[13119:13112];
        434: state_byte <= hashes[13111:13104];
        435: state_byte <= hashes[13103:13096];
        436: state_byte <= hashes[13095:13088];
        437: state_byte <= hashes[13087:13080];
        438: state_byte <= hashes[13079:13072];
        439: state_byte <= hashes[13071:13064];
        440: state_byte <= hashes[13063:13056];
        441: state_byte <= hashes[13055:13048];
        442: state_byte <= hashes[13047:13040];
        443: state_byte <= hashes[13039:13032];
        444: state_byte <= hashes[13031:13024];
        445: state_byte <= hashes[13023:13016];
        446: state_byte <= hashes[13015:13008];
        447: state_byte <= hashes[13007:13000];
        448: state_byte <= hashes[12999:12992];
        449: state_byte <= hashes[12991:12984];
        450: state_byte <= hashes[12983:12976];
        451: state_byte <= hashes[12975:12968];
        452: state_byte <= hashes[12967:12960];
        453: state_byte <= hashes[12959:12952];
        454: state_byte <= hashes[12951:12944];
        455: state_byte <= hashes[12943:12936];
        456: state_byte <= hashes[12935:12928];
        457: state_byte <= hashes[12927:12920];
        458: state_byte <= hashes[12919:12912];
        459: state_byte <= hashes[12911:12904];
        460: state_byte <= hashes[12903:12896];
        461: state_byte <= hashes[12895:12888];
        462: state_byte <= hashes[12887:12880];
        463: state_byte <= hashes[12879:12872];
        464: state_byte <= hashes[12871:12864];
        465: state_byte <= hashes[12863:12856];
        466: state_byte <= hashes[12855:12848];
        467: state_byte <= hashes[12847:12840];
        468: state_byte <= hashes[12839:12832];
        469: state_byte <= hashes[12831:12824];
        470: state_byte <= hashes[12823:12816];
        471: state_byte <= hashes[12815:12808];
        472: state_byte <= hashes[12807:12800];
        473: state_byte <= hashes[12799:12792];
        474: state_byte <= hashes[12791:12784];
        475: state_byte <= hashes[12783:12776];
        476: state_byte <= hashes[12775:12768];
        477: state_byte <= hashes[12767:12760];
        478: state_byte <= hashes[12759:12752];
        479: state_byte <= hashes[12751:12744];
        480: state_byte <= hashes[12743:12736];
        481: state_byte <= hashes[12735:12728];
        482: state_byte <= hashes[12727:12720];
        483: state_byte <= hashes[12719:12712];
        484: state_byte <= hashes[12711:12704];
        485: state_byte <= hashes[12703:12696];
        486: state_byte <= hashes[12695:12688];
        487: state_byte <= hashes[12687:12680];
        488: state_byte <= hashes[12679:12672];
        489: state_byte <= hashes[12671:12664];
        490: state_byte <= hashes[12663:12656];
        491: state_byte <= hashes[12655:12648];
        492: state_byte <= hashes[12647:12640];
        493: state_byte <= hashes[12639:12632];
        494: state_byte <= hashes[12631:12624];
        495: state_byte <= hashes[12623:12616];
        496: state_byte <= hashes[12615:12608];
        497: state_byte <= hashes[12607:12600];
        498: state_byte <= hashes[12599:12592];
        499: state_byte <= hashes[12591:12584];
        500: state_byte <= hashes[12583:12576];
        501: state_byte <= hashes[12575:12568];
        502: state_byte <= hashes[12567:12560];
        503: state_byte <= hashes[12559:12552];
        504: state_byte <= hashes[12551:12544];
        505: state_byte <= hashes[12543:12536];
        506: state_byte <= hashes[12535:12528];
        507: state_byte <= hashes[12527:12520];
        508: state_byte <= hashes[12519:12512];
        509: state_byte <= hashes[12511:12504];
        510: state_byte <= hashes[12503:12496];
        511: state_byte <= hashes[12495:12488];
        512: state_byte <= hashes[12487:12480];
        513: state_byte <= hashes[12479:12472];
        514: state_byte <= hashes[12471:12464];
        515: state_byte <= hashes[12463:12456];
        516: state_byte <= hashes[12455:12448];
        517: state_byte <= hashes[12447:12440];
        518: state_byte <= hashes[12439:12432];
        519: state_byte <= hashes[12431:12424];
        520: state_byte <= hashes[12423:12416];
        521: state_byte <= hashes[12415:12408];
        522: state_byte <= hashes[12407:12400];
        523: state_byte <= hashes[12399:12392];
        524: state_byte <= hashes[12391:12384];
        525: state_byte <= hashes[12383:12376];
        526: state_byte <= hashes[12375:12368];
        527: state_byte <= hashes[12367:12360];
        528: state_byte <= hashes[12359:12352];
        529: state_byte <= hashes[12351:12344];
        530: state_byte <= hashes[12343:12336];
        531: state_byte <= hashes[12335:12328];
        532: state_byte <= hashes[12327:12320];
        533: state_byte <= hashes[12319:12312];
        534: state_byte <= hashes[12311:12304];
        535: state_byte <= hashes[12303:12296];
        536: state_byte <= hashes[12295:12288];
        537: state_byte <= hashes[12287:12280];
        538: state_byte <= hashes[12279:12272];
        539: state_byte <= hashes[12271:12264];
        540: state_byte <= hashes[12263:12256];
        541: state_byte <= hashes[12255:12248];
        542: state_byte <= hashes[12247:12240];
        543: state_byte <= hashes[12239:12232];
        544: state_byte <= hashes[12231:12224];
        545: state_byte <= hashes[12223:12216];
        546: state_byte <= hashes[12215:12208];
        547: state_byte <= hashes[12207:12200];
        548: state_byte <= hashes[12199:12192];
        549: state_byte <= hashes[12191:12184];
        550: state_byte <= hashes[12183:12176];
        551: state_byte <= hashes[12175:12168];
        552: state_byte <= hashes[12167:12160];
        553: state_byte <= hashes[12159:12152];
        554: state_byte <= hashes[12151:12144];
        555: state_byte <= hashes[12143:12136];
        556: state_byte <= hashes[12135:12128];
        557: state_byte <= hashes[12127:12120];
        558: state_byte <= hashes[12119:12112];
        559: state_byte <= hashes[12111:12104];
        560: state_byte <= hashes[12103:12096];
        561: state_byte <= hashes[12095:12088];
        562: state_byte <= hashes[12087:12080];
        563: state_byte <= hashes[12079:12072];
        564: state_byte <= hashes[12071:12064];
        565: state_byte <= hashes[12063:12056];
        566: state_byte <= hashes[12055:12048];
        567: state_byte <= hashes[12047:12040];
        568: state_byte <= hashes[12039:12032];
        569: state_byte <= hashes[12031:12024];
        570: state_byte <= hashes[12023:12016];
        571: state_byte <= hashes[12015:12008];
        572: state_byte <= hashes[12007:12000];
        573: state_byte <= hashes[11999:11992];
        574: state_byte <= hashes[11991:11984];
        575: state_byte <= hashes[11983:11976];
        576: state_byte <= hashes[11975:11968];
        577: state_byte <= hashes[11967:11960];
        578: state_byte <= hashes[11959:11952];
        579: state_byte <= hashes[11951:11944];
        580: state_byte <= hashes[11943:11936];
        581: state_byte <= hashes[11935:11928];
        582: state_byte <= hashes[11927:11920];
        583: state_byte <= hashes[11919:11912];
        584: state_byte <= hashes[11911:11904];
        585: state_byte <= hashes[11903:11896];
        586: state_byte <= hashes[11895:11888];
        587: state_byte <= hashes[11887:11880];
        588: state_byte <= hashes[11879:11872];
        589: state_byte <= hashes[11871:11864];
        590: state_byte <= hashes[11863:11856];
        591: state_byte <= hashes[11855:11848];
        592: state_byte <= hashes[11847:11840];
        593: state_byte <= hashes[11839:11832];
        594: state_byte <= hashes[11831:11824];
        595: state_byte <= hashes[11823:11816];
        596: state_byte <= hashes[11815:11808];
        597: state_byte <= hashes[11807:11800];
        598: state_byte <= hashes[11799:11792];
        599: state_byte <= hashes[11791:11784];
        600: state_byte <= hashes[11783:11776];
        601: state_byte <= hashes[11775:11768];
        602: state_byte <= hashes[11767:11760];
        603: state_byte <= hashes[11759:11752];
        604: state_byte <= hashes[11751:11744];
        605: state_byte <= hashes[11743:11736];
        606: state_byte <= hashes[11735:11728];
        607: state_byte <= hashes[11727:11720];
        608: state_byte <= hashes[11719:11712];
        609: state_byte <= hashes[11711:11704];
        610: state_byte <= hashes[11703:11696];
        611: state_byte <= hashes[11695:11688];
        612: state_byte <= hashes[11687:11680];
        613: state_byte <= hashes[11679:11672];
        614: state_byte <= hashes[11671:11664];
        615: state_byte <= hashes[11663:11656];
        616: state_byte <= hashes[11655:11648];
        617: state_byte <= hashes[11647:11640];
        618: state_byte <= hashes[11639:11632];
        619: state_byte <= hashes[11631:11624];
        620: state_byte <= hashes[11623:11616];
        621: state_byte <= hashes[11615:11608];
        622: state_byte <= hashes[11607:11600];
        623: state_byte <= hashes[11599:11592];
        624: state_byte <= hashes[11591:11584];
        625: state_byte <= hashes[11583:11576];
        626: state_byte <= hashes[11575:11568];
        627: state_byte <= hashes[11567:11560];
        628: state_byte <= hashes[11559:11552];
        629: state_byte <= hashes[11551:11544];
        630: state_byte <= hashes[11543:11536];
        631: state_byte <= hashes[11535:11528];
        632: state_byte <= hashes[11527:11520];
        633: state_byte <= hashes[11519:11512];
        634: state_byte <= hashes[11511:11504];
        635: state_byte <= hashes[11503:11496];
        636: state_byte <= hashes[11495:11488];
        637: state_byte <= hashes[11487:11480];
        638: state_byte <= hashes[11479:11472];
        639: state_byte <= hashes[11471:11464];
        640: state_byte <= hashes[11463:11456];
        641: state_byte <= hashes[11455:11448];
        642: state_byte <= hashes[11447:11440];
        643: state_byte <= hashes[11439:11432];
        644: state_byte <= hashes[11431:11424];
        645: state_byte <= hashes[11423:11416];
        646: state_byte <= hashes[11415:11408];
        647: state_byte <= hashes[11407:11400];
        648: state_byte <= hashes[11399:11392];
        649: state_byte <= hashes[11391:11384];
        650: state_byte <= hashes[11383:11376];
        651: state_byte <= hashes[11375:11368];
        652: state_byte <= hashes[11367:11360];
        653: state_byte <= hashes[11359:11352];
        654: state_byte <= hashes[11351:11344];
        655: state_byte <= hashes[11343:11336];
        656: state_byte <= hashes[11335:11328];
        657: state_byte <= hashes[11327:11320];
        658: state_byte <= hashes[11319:11312];
        659: state_byte <= hashes[11311:11304];
        660: state_byte <= hashes[11303:11296];
        661: state_byte <= hashes[11295:11288];
        662: state_byte <= hashes[11287:11280];
        663: state_byte <= hashes[11279:11272];
        664: state_byte <= hashes[11271:11264];
        665: state_byte <= hashes[11263:11256];
        666: state_byte <= hashes[11255:11248];
        667: state_byte <= hashes[11247:11240];
        668: state_byte <= hashes[11239:11232];
        669: state_byte <= hashes[11231:11224];
        670: state_byte <= hashes[11223:11216];
        671: state_byte <= hashes[11215:11208];
        672: state_byte <= hashes[11207:11200];
        673: state_byte <= hashes[11199:11192];
        674: state_byte <= hashes[11191:11184];
        675: state_byte <= hashes[11183:11176];
        676: state_byte <= hashes[11175:11168];
        677: state_byte <= hashes[11167:11160];
        678: state_byte <= hashes[11159:11152];
        679: state_byte <= hashes[11151:11144];
        680: state_byte <= hashes[11143:11136];
        681: state_byte <= hashes[11135:11128];
        682: state_byte <= hashes[11127:11120];
        683: state_byte <= hashes[11119:11112];
        684: state_byte <= hashes[11111:11104];
        685: state_byte <= hashes[11103:11096];
        686: state_byte <= hashes[11095:11088];
        687: state_byte <= hashes[11087:11080];
        688: state_byte <= hashes[11079:11072];
        689: state_byte <= hashes[11071:11064];
        690: state_byte <= hashes[11063:11056];
        691: state_byte <= hashes[11055:11048];
        692: state_byte <= hashes[11047:11040];
        693: state_byte <= hashes[11039:11032];
        694: state_byte <= hashes[11031:11024];
        695: state_byte <= hashes[11023:11016];
        696: state_byte <= hashes[11015:11008];
        697: state_byte <= hashes[11007:11000];
        698: state_byte <= hashes[10999:10992];
        699: state_byte <= hashes[10991:10984];
        700: state_byte <= hashes[10983:10976];
        701: state_byte <= hashes[10975:10968];
        702: state_byte <= hashes[10967:10960];
        703: state_byte <= hashes[10959:10952];
        704: state_byte <= hashes[10951:10944];
        705: state_byte <= hashes[10943:10936];
        706: state_byte <= hashes[10935:10928];
        707: state_byte <= hashes[10927:10920];
        708: state_byte <= hashes[10919:10912];
        709: state_byte <= hashes[10911:10904];
        710: state_byte <= hashes[10903:10896];
        711: state_byte <= hashes[10895:10888];
        712: state_byte <= hashes[10887:10880];
        713: state_byte <= hashes[10879:10872];
        714: state_byte <= hashes[10871:10864];
        715: state_byte <= hashes[10863:10856];
        716: state_byte <= hashes[10855:10848];
        717: state_byte <= hashes[10847:10840];
        718: state_byte <= hashes[10839:10832];
        719: state_byte <= hashes[10831:10824];
        720: state_byte <= hashes[10823:10816];
        721: state_byte <= hashes[10815:10808];
        722: state_byte <= hashes[10807:10800];
        723: state_byte <= hashes[10799:10792];
        724: state_byte <= hashes[10791:10784];
        725: state_byte <= hashes[10783:10776];
        726: state_byte <= hashes[10775:10768];
        727: state_byte <= hashes[10767:10760];
        728: state_byte <= hashes[10759:10752];
        729: state_byte <= hashes[10751:10744];
        730: state_byte <= hashes[10743:10736];
        731: state_byte <= hashes[10735:10728];
        732: state_byte <= hashes[10727:10720];
        733: state_byte <= hashes[10719:10712];
        734: state_byte <= hashes[10711:10704];
        735: state_byte <= hashes[10703:10696];
        736: state_byte <= hashes[10695:10688];
        737: state_byte <= hashes[10687:10680];
        738: state_byte <= hashes[10679:10672];
        739: state_byte <= hashes[10671:10664];
        740: state_byte <= hashes[10663:10656];
        741: state_byte <= hashes[10655:10648];
        742: state_byte <= hashes[10647:10640];
        743: state_byte <= hashes[10639:10632];
        744: state_byte <= hashes[10631:10624];
        745: state_byte <= hashes[10623:10616];
        746: state_byte <= hashes[10615:10608];
        747: state_byte <= hashes[10607:10600];
        748: state_byte <= hashes[10599:10592];
        749: state_byte <= hashes[10591:10584];
        750: state_byte <= hashes[10583:10576];
        751: state_byte <= hashes[10575:10568];
        752: state_byte <= hashes[10567:10560];
        753: state_byte <= hashes[10559:10552];
        754: state_byte <= hashes[10551:10544];
        755: state_byte <= hashes[10543:10536];
        756: state_byte <= hashes[10535:10528];
        757: state_byte <= hashes[10527:10520];
        758: state_byte <= hashes[10519:10512];
        759: state_byte <= hashes[10511:10504];
        760: state_byte <= hashes[10503:10496];
        761: state_byte <= hashes[10495:10488];
        762: state_byte <= hashes[10487:10480];
        763: state_byte <= hashes[10479:10472];
        764: state_byte <= hashes[10471:10464];
        765: state_byte <= hashes[10463:10456];
        766: state_byte <= hashes[10455:10448];
        767: state_byte <= hashes[10447:10440];
        768: state_byte <= hashes[10439:10432];
        769: state_byte <= hashes[10431:10424];
        770: state_byte <= hashes[10423:10416];
        771: state_byte <= hashes[10415:10408];
        772: state_byte <= hashes[10407:10400];
        773: state_byte <= hashes[10399:10392];
        774: state_byte <= hashes[10391:10384];
        775: state_byte <= hashes[10383:10376];
        776: state_byte <= hashes[10375:10368];
        777: state_byte <= hashes[10367:10360];
        778: state_byte <= hashes[10359:10352];
        779: state_byte <= hashes[10351:10344];
        780: state_byte <= hashes[10343:10336];
        781: state_byte <= hashes[10335:10328];
        782: state_byte <= hashes[10327:10320];
        783: state_byte <= hashes[10319:10312];
        784: state_byte <= hashes[10311:10304];
        785: state_byte <= hashes[10303:10296];
        786: state_byte <= hashes[10295:10288];
        787: state_byte <= hashes[10287:10280];
        788: state_byte <= hashes[10279:10272];
        789: state_byte <= hashes[10271:10264];
        790: state_byte <= hashes[10263:10256];
        791: state_byte <= hashes[10255:10248];
        792: state_byte <= hashes[10247:10240];
        793: state_byte <= hashes[10239:10232];
        794: state_byte <= hashes[10231:10224];
        795: state_byte <= hashes[10223:10216];
        796: state_byte <= hashes[10215:10208];
        797: state_byte <= hashes[10207:10200];
        798: state_byte <= hashes[10199:10192];
        799: state_byte <= hashes[10191:10184];
        800: state_byte <= hashes[10183:10176];
        801: state_byte <= hashes[10175:10168];
        802: state_byte <= hashes[10167:10160];
        803: state_byte <= hashes[10159:10152];
        804: state_byte <= hashes[10151:10144];
        805: state_byte <= hashes[10143:10136];
        806: state_byte <= hashes[10135:10128];
        807: state_byte <= hashes[10127:10120];
        808: state_byte <= hashes[10119:10112];
        809: state_byte <= hashes[10111:10104];
        810: state_byte <= hashes[10103:10096];
        811: state_byte <= hashes[10095:10088];
        812: state_byte <= hashes[10087:10080];
        813: state_byte <= hashes[10079:10072];
        814: state_byte <= hashes[10071:10064];
        815: state_byte <= hashes[10063:10056];
        816: state_byte <= hashes[10055:10048];
        817: state_byte <= hashes[10047:10040];
        818: state_byte <= hashes[10039:10032];
        819: state_byte <= hashes[10031:10024];
        820: state_byte <= hashes[10023:10016];
        821: state_byte <= hashes[10015:10008];
        822: state_byte <= hashes[10007:10000];
        823: state_byte <= hashes[9999:9992];
        824: state_byte <= hashes[9991:9984];
        825: state_byte <= hashes[9983:9976];
        826: state_byte <= hashes[9975:9968];
        827: state_byte <= hashes[9967:9960];
        828: state_byte <= hashes[9959:9952];
        829: state_byte <= hashes[9951:9944];
        830: state_byte <= hashes[9943:9936];
        831: state_byte <= hashes[9935:9928];
        832: state_byte <= hashes[9927:9920];
        833: state_byte <= hashes[9919:9912];
        834: state_byte <= hashes[9911:9904];
        835: state_byte <= hashes[9903:9896];
        836: state_byte <= hashes[9895:9888];
        837: state_byte <= hashes[9887:9880];
        838: state_byte <= hashes[9879:9872];
        839: state_byte <= hashes[9871:9864];
        840: state_byte <= hashes[9863:9856];
        841: state_byte <= hashes[9855:9848];
        842: state_byte <= hashes[9847:9840];
        843: state_byte <= hashes[9839:9832];
        844: state_byte <= hashes[9831:9824];
        845: state_byte <= hashes[9823:9816];
        846: state_byte <= hashes[9815:9808];
        847: state_byte <= hashes[9807:9800];
        848: state_byte <= hashes[9799:9792];
        849: state_byte <= hashes[9791:9784];
        850: state_byte <= hashes[9783:9776];
        851: state_byte <= hashes[9775:9768];
        852: state_byte <= hashes[9767:9760];
        853: state_byte <= hashes[9759:9752];
        854: state_byte <= hashes[9751:9744];
        855: state_byte <= hashes[9743:9736];
        856: state_byte <= hashes[9735:9728];
        857: state_byte <= hashes[9727:9720];
        858: state_byte <= hashes[9719:9712];
        859: state_byte <= hashes[9711:9704];
        860: state_byte <= hashes[9703:9696];
        861: state_byte <= hashes[9695:9688];
        862: state_byte <= hashes[9687:9680];
        863: state_byte <= hashes[9679:9672];
        864: state_byte <= hashes[9671:9664];
        865: state_byte <= hashes[9663:9656];
        866: state_byte <= hashes[9655:9648];
        867: state_byte <= hashes[9647:9640];
        868: state_byte <= hashes[9639:9632];
        869: state_byte <= hashes[9631:9624];
        870: state_byte <= hashes[9623:9616];
        871: state_byte <= hashes[9615:9608];
        872: state_byte <= hashes[9607:9600];
        873: state_byte <= hashes[9599:9592];
        874: state_byte <= hashes[9591:9584];
        875: state_byte <= hashes[9583:9576];
        876: state_byte <= hashes[9575:9568];
        877: state_byte <= hashes[9567:9560];
        878: state_byte <= hashes[9559:9552];
        879: state_byte <= hashes[9551:9544];
        880: state_byte <= hashes[9543:9536];
        881: state_byte <= hashes[9535:9528];
        882: state_byte <= hashes[9527:9520];
        883: state_byte <= hashes[9519:9512];
        884: state_byte <= hashes[9511:9504];
        885: state_byte <= hashes[9503:9496];
        886: state_byte <= hashes[9495:9488];
        887: state_byte <= hashes[9487:9480];
        888: state_byte <= hashes[9479:9472];
        889: state_byte <= hashes[9471:9464];
        890: state_byte <= hashes[9463:9456];
        891: state_byte <= hashes[9455:9448];
        892: state_byte <= hashes[9447:9440];
        893: state_byte <= hashes[9439:9432];
        894: state_byte <= hashes[9431:9424];
        895: state_byte <= hashes[9423:9416];
        896: state_byte <= hashes[9415:9408];
        897: state_byte <= hashes[9407:9400];
        898: state_byte <= hashes[9399:9392];
        899: state_byte <= hashes[9391:9384];
        900: state_byte <= hashes[9383:9376];
        901: state_byte <= hashes[9375:9368];
        902: state_byte <= hashes[9367:9360];
        903: state_byte <= hashes[9359:9352];
        904: state_byte <= hashes[9351:9344];
        905: state_byte <= hashes[9343:9336];
        906: state_byte <= hashes[9335:9328];
        907: state_byte <= hashes[9327:9320];
        908: state_byte <= hashes[9319:9312];
        909: state_byte <= hashes[9311:9304];
        910: state_byte <= hashes[9303:9296];
        911: state_byte <= hashes[9295:9288];
        912: state_byte <= hashes[9287:9280];
        913: state_byte <= hashes[9279:9272];
        914: state_byte <= hashes[9271:9264];
        915: state_byte <= hashes[9263:9256];
        916: state_byte <= hashes[9255:9248];
        917: state_byte <= hashes[9247:9240];
        918: state_byte <= hashes[9239:9232];
        919: state_byte <= hashes[9231:9224];
        920: state_byte <= hashes[9223:9216];
        921: state_byte <= hashes[9215:9208];
        922: state_byte <= hashes[9207:9200];
        923: state_byte <= hashes[9199:9192];
        924: state_byte <= hashes[9191:9184];
        925: state_byte <= hashes[9183:9176];
        926: state_byte <= hashes[9175:9168];
        927: state_byte <= hashes[9167:9160];
        928: state_byte <= hashes[9159:9152];
        929: state_byte <= hashes[9151:9144];
        930: state_byte <= hashes[9143:9136];
        931: state_byte <= hashes[9135:9128];
        932: state_byte <= hashes[9127:9120];
        933: state_byte <= hashes[9119:9112];
        934: state_byte <= hashes[9111:9104];
        935: state_byte <= hashes[9103:9096];
        936: state_byte <= hashes[9095:9088];
        937: state_byte <= hashes[9087:9080];
        938: state_byte <= hashes[9079:9072];
        939: state_byte <= hashes[9071:9064];
        940: state_byte <= hashes[9063:9056];
        941: state_byte <= hashes[9055:9048];
        942: state_byte <= hashes[9047:9040];
        943: state_byte <= hashes[9039:9032];
        944: state_byte <= hashes[9031:9024];
        945: state_byte <= hashes[9023:9016];
        946: state_byte <= hashes[9015:9008];
        947: state_byte <= hashes[9007:9000];
        948: state_byte <= hashes[8999:8992];
        949: state_byte <= hashes[8991:8984];
        950: state_byte <= hashes[8983:8976];
        951: state_byte <= hashes[8975:8968];
        952: state_byte <= hashes[8967:8960];
        953: state_byte <= hashes[8959:8952];
        954: state_byte <= hashes[8951:8944];
        955: state_byte <= hashes[8943:8936];
        956: state_byte <= hashes[8935:8928];
        957: state_byte <= hashes[8927:8920];
        958: state_byte <= hashes[8919:8912];
        959: state_byte <= hashes[8911:8904];
        960: state_byte <= hashes[8903:8896];
        961: state_byte <= hashes[8895:8888];
        962: state_byte <= hashes[8887:8880];
        963: state_byte <= hashes[8879:8872];
        964: state_byte <= hashes[8871:8864];
        965: state_byte <= hashes[8863:8856];
        966: state_byte <= hashes[8855:8848];
        967: state_byte <= hashes[8847:8840];
        968: state_byte <= hashes[8839:8832];
        969: state_byte <= hashes[8831:8824];
        970: state_byte <= hashes[8823:8816];
        971: state_byte <= hashes[8815:8808];
        972: state_byte <= hashes[8807:8800];
        973: state_byte <= hashes[8799:8792];
        974: state_byte <= hashes[8791:8784];
        975: state_byte <= hashes[8783:8776];
        976: state_byte <= hashes[8775:8768];
        977: state_byte <= hashes[8767:8760];
        978: state_byte <= hashes[8759:8752];
        979: state_byte <= hashes[8751:8744];
        980: state_byte <= hashes[8743:8736];
        981: state_byte <= hashes[8735:8728];
        982: state_byte <= hashes[8727:8720];
        983: state_byte <= hashes[8719:8712];
        984: state_byte <= hashes[8711:8704];
        985: state_byte <= hashes[8703:8696];
        986: state_byte <= hashes[8695:8688];
        987: state_byte <= hashes[8687:8680];
        988: state_byte <= hashes[8679:8672];
        989: state_byte <= hashes[8671:8664];
        990: state_byte <= hashes[8663:8656];
        991: state_byte <= hashes[8655:8648];
        992: state_byte <= hashes[8647:8640];
        993: state_byte <= hashes[8639:8632];
        994: state_byte <= hashes[8631:8624];
        995: state_byte <= hashes[8623:8616];
        996: state_byte <= hashes[8615:8608];
        997: state_byte <= hashes[8607:8600];
        998: state_byte <= hashes[8599:8592];
        999: state_byte <= hashes[8591:8584];
        1000: state_byte <= hashes[8583:8576];
        1001: state_byte <= hashes[8575:8568];
        1002: state_byte <= hashes[8567:8560];
        1003: state_byte <= hashes[8559:8552];
        1004: state_byte <= hashes[8551:8544];
        1005: state_byte <= hashes[8543:8536];
        1006: state_byte <= hashes[8535:8528];
        1007: state_byte <= hashes[8527:8520];
        1008: state_byte <= hashes[8519:8512];
        1009: state_byte <= hashes[8511:8504];
        1010: state_byte <= hashes[8503:8496];
        1011: state_byte <= hashes[8495:8488];
        1012: state_byte <= hashes[8487:8480];
        1013: state_byte <= hashes[8479:8472];
        1014: state_byte <= hashes[8471:8464];
        1015: state_byte <= hashes[8463:8456];
        1016: state_byte <= hashes[8455:8448];
        1017: state_byte <= hashes[8447:8440];
        1018: state_byte <= hashes[8439:8432];
        1019: state_byte <= hashes[8431:8424];
        1020: state_byte <= hashes[8423:8416];
        1021: state_byte <= hashes[8415:8408];
        1022: state_byte <= hashes[8407:8400];
        1023: state_byte <= hashes[8399:8392];
        1024: state_byte <= hashes[8391:8384];
        1025: state_byte <= hashes[8383:8376];
        1026: state_byte <= hashes[8375:8368];
        1027: state_byte <= hashes[8367:8360];
        1028: state_byte <= hashes[8359:8352];
        1029: state_byte <= hashes[8351:8344];
        1030: state_byte <= hashes[8343:8336];
        1031: state_byte <= hashes[8335:8328];
        1032: state_byte <= hashes[8327:8320];
        1033: state_byte <= hashes[8319:8312];
        1034: state_byte <= hashes[8311:8304];
        1035: state_byte <= hashes[8303:8296];
        1036: state_byte <= hashes[8295:8288];
        1037: state_byte <= hashes[8287:8280];
        1038: state_byte <= hashes[8279:8272];
        1039: state_byte <= hashes[8271:8264];
        1040: state_byte <= hashes[8263:8256];
        1041: state_byte <= hashes[8255:8248];
        1042: state_byte <= hashes[8247:8240];
        1043: state_byte <= hashes[8239:8232];
        1044: state_byte <= hashes[8231:8224];
        1045: state_byte <= hashes[8223:8216];
        1046: state_byte <= hashes[8215:8208];
        1047: state_byte <= hashes[8207:8200];
        1048: state_byte <= hashes[8199:8192];
        1049: state_byte <= hashes[8191:8184];
        1050: state_byte <= hashes[8183:8176];
        1051: state_byte <= hashes[8175:8168];
        1052: state_byte <= hashes[8167:8160];
        1053: state_byte <= hashes[8159:8152];
        1054: state_byte <= hashes[8151:8144];
        1055: state_byte <= hashes[8143:8136];
        1056: state_byte <= hashes[8135:8128];
        1057: state_byte <= hashes[8127:8120];
        1058: state_byte <= hashes[8119:8112];
        1059: state_byte <= hashes[8111:8104];
        1060: state_byte <= hashes[8103:8096];
        1061: state_byte <= hashes[8095:8088];
        1062: state_byte <= hashes[8087:8080];
        1063: state_byte <= hashes[8079:8072];
        1064: state_byte <= hashes[8071:8064];
        1065: state_byte <= hashes[8063:8056];
        1066: state_byte <= hashes[8055:8048];
        1067: state_byte <= hashes[8047:8040];
        1068: state_byte <= hashes[8039:8032];
        1069: state_byte <= hashes[8031:8024];
        1070: state_byte <= hashes[8023:8016];
        1071: state_byte <= hashes[8015:8008];
        1072: state_byte <= hashes[8007:8000];
        1073: state_byte <= hashes[7999:7992];
        1074: state_byte <= hashes[7991:7984];
        1075: state_byte <= hashes[7983:7976];
        1076: state_byte <= hashes[7975:7968];
        1077: state_byte <= hashes[7967:7960];
        1078: state_byte <= hashes[7959:7952];
        1079: state_byte <= hashes[7951:7944];
        1080: state_byte <= hashes[7943:7936];
        1081: state_byte <= hashes[7935:7928];
        1082: state_byte <= hashes[7927:7920];
        1083: state_byte <= hashes[7919:7912];
        1084: state_byte <= hashes[7911:7904];
        1085: state_byte <= hashes[7903:7896];
        1086: state_byte <= hashes[7895:7888];
        1087: state_byte <= hashes[7887:7880];
        1088: state_byte <= hashes[7879:7872];
        1089: state_byte <= hashes[7871:7864];
        1090: state_byte <= hashes[7863:7856];
        1091: state_byte <= hashes[7855:7848];
        1092: state_byte <= hashes[7847:7840];
        1093: state_byte <= hashes[7839:7832];
        1094: state_byte <= hashes[7831:7824];
        1095: state_byte <= hashes[7823:7816];
        1096: state_byte <= hashes[7815:7808];
        1097: state_byte <= hashes[7807:7800];
        1098: state_byte <= hashes[7799:7792];
        1099: state_byte <= hashes[7791:7784];
        1100: state_byte <= hashes[7783:7776];
        1101: state_byte <= hashes[7775:7768];
        1102: state_byte <= hashes[7767:7760];
        1103: state_byte <= hashes[7759:7752];
        1104: state_byte <= hashes[7751:7744];
        1105: state_byte <= hashes[7743:7736];
        1106: state_byte <= hashes[7735:7728];
        1107: state_byte <= hashes[7727:7720];
        1108: state_byte <= hashes[7719:7712];
        1109: state_byte <= hashes[7711:7704];
        1110: state_byte <= hashes[7703:7696];
        1111: state_byte <= hashes[7695:7688];
        1112: state_byte <= hashes[7687:7680];
        1113: state_byte <= hashes[7679:7672];
        1114: state_byte <= hashes[7671:7664];
        1115: state_byte <= hashes[7663:7656];
        1116: state_byte <= hashes[7655:7648];
        1117: state_byte <= hashes[7647:7640];
        1118: state_byte <= hashes[7639:7632];
        1119: state_byte <= hashes[7631:7624];
        1120: state_byte <= hashes[7623:7616];
        1121: state_byte <= hashes[7615:7608];
        1122: state_byte <= hashes[7607:7600];
        1123: state_byte <= hashes[7599:7592];
        1124: state_byte <= hashes[7591:7584];
        1125: state_byte <= hashes[7583:7576];
        1126: state_byte <= hashes[7575:7568];
        1127: state_byte <= hashes[7567:7560];
        1128: state_byte <= hashes[7559:7552];
        1129: state_byte <= hashes[7551:7544];
        1130: state_byte <= hashes[7543:7536];
        1131: state_byte <= hashes[7535:7528];
        1132: state_byte <= hashes[7527:7520];
        1133: state_byte <= hashes[7519:7512];
        1134: state_byte <= hashes[7511:7504];
        1135: state_byte <= hashes[7503:7496];
        1136: state_byte <= hashes[7495:7488];
        1137: state_byte <= hashes[7487:7480];
        1138: state_byte <= hashes[7479:7472];
        1139: state_byte <= hashes[7471:7464];
        1140: state_byte <= hashes[7463:7456];
        1141: state_byte <= hashes[7455:7448];
        1142: state_byte <= hashes[7447:7440];
        1143: state_byte <= hashes[7439:7432];
        1144: state_byte <= hashes[7431:7424];
        1145: state_byte <= hashes[7423:7416];
        1146: state_byte <= hashes[7415:7408];
        1147: state_byte <= hashes[7407:7400];
        1148: state_byte <= hashes[7399:7392];
        1149: state_byte <= hashes[7391:7384];
        1150: state_byte <= hashes[7383:7376];
        1151: state_byte <= hashes[7375:7368];
        1152: state_byte <= hashes[7367:7360];
        1153: state_byte <= hashes[7359:7352];
        1154: state_byte <= hashes[7351:7344];
        1155: state_byte <= hashes[7343:7336];
        1156: state_byte <= hashes[7335:7328];
        1157: state_byte <= hashes[7327:7320];
        1158: state_byte <= hashes[7319:7312];
        1159: state_byte <= hashes[7311:7304];
        1160: state_byte <= hashes[7303:7296];
        1161: state_byte <= hashes[7295:7288];
        1162: state_byte <= hashes[7287:7280];
        1163: state_byte <= hashes[7279:7272];
        1164: state_byte <= hashes[7271:7264];
        1165: state_byte <= hashes[7263:7256];
        1166: state_byte <= hashes[7255:7248];
        1167: state_byte <= hashes[7247:7240];
        1168: state_byte <= hashes[7239:7232];
        1169: state_byte <= hashes[7231:7224];
        1170: state_byte <= hashes[7223:7216];
        1171: state_byte <= hashes[7215:7208];
        1172: state_byte <= hashes[7207:7200];
        1173: state_byte <= hashes[7199:7192];
        1174: state_byte <= hashes[7191:7184];
        1175: state_byte <= hashes[7183:7176];
        1176: state_byte <= hashes[7175:7168];
        1177: state_byte <= hashes[7167:7160];
        1178: state_byte <= hashes[7159:7152];
        1179: state_byte <= hashes[7151:7144];
        1180: state_byte <= hashes[7143:7136];
        1181: state_byte <= hashes[7135:7128];
        1182: state_byte <= hashes[7127:7120];
        1183: state_byte <= hashes[7119:7112];
        1184: state_byte <= hashes[7111:7104];
        1185: state_byte <= hashes[7103:7096];
        1186: state_byte <= hashes[7095:7088];
        1187: state_byte <= hashes[7087:7080];
        1188: state_byte <= hashes[7079:7072];
        1189: state_byte <= hashes[7071:7064];
        1190: state_byte <= hashes[7063:7056];
        1191: state_byte <= hashes[7055:7048];
        1192: state_byte <= hashes[7047:7040];
        1193: state_byte <= hashes[7039:7032];
        1194: state_byte <= hashes[7031:7024];
        1195: state_byte <= hashes[7023:7016];
        1196: state_byte <= hashes[7015:7008];
        1197: state_byte <= hashes[7007:7000];
        1198: state_byte <= hashes[6999:6992];
        1199: state_byte <= hashes[6991:6984];
        1200: state_byte <= hashes[6983:6976];
        1201: state_byte <= hashes[6975:6968];
        1202: state_byte <= hashes[6967:6960];
        1203: state_byte <= hashes[6959:6952];
        1204: state_byte <= hashes[6951:6944];
        1205: state_byte <= hashes[6943:6936];
        1206: state_byte <= hashes[6935:6928];
        1207: state_byte <= hashes[6927:6920];
        1208: state_byte <= hashes[6919:6912];
        1209: state_byte <= hashes[6911:6904];
        1210: state_byte <= hashes[6903:6896];
        1211: state_byte <= hashes[6895:6888];
        1212: state_byte <= hashes[6887:6880];
        1213: state_byte <= hashes[6879:6872];
        1214: state_byte <= hashes[6871:6864];
        1215: state_byte <= hashes[6863:6856];
        1216: state_byte <= hashes[6855:6848];
        1217: state_byte <= hashes[6847:6840];
        1218: state_byte <= hashes[6839:6832];
        1219: state_byte <= hashes[6831:6824];
        1220: state_byte <= hashes[6823:6816];
        1221: state_byte <= hashes[6815:6808];
        1222: state_byte <= hashes[6807:6800];
        1223: state_byte <= hashes[6799:6792];
        1224: state_byte <= hashes[6791:6784];
        1225: state_byte <= hashes[6783:6776];
        1226: state_byte <= hashes[6775:6768];
        1227: state_byte <= hashes[6767:6760];
        1228: state_byte <= hashes[6759:6752];
        1229: state_byte <= hashes[6751:6744];
        1230: state_byte <= hashes[6743:6736];
        1231: state_byte <= hashes[6735:6728];
        1232: state_byte <= hashes[6727:6720];
        1233: state_byte <= hashes[6719:6712];
        1234: state_byte <= hashes[6711:6704];
        1235: state_byte <= hashes[6703:6696];
        1236: state_byte <= hashes[6695:6688];
        1237: state_byte <= hashes[6687:6680];
        1238: state_byte <= hashes[6679:6672];
        1239: state_byte <= hashes[6671:6664];
        1240: state_byte <= hashes[6663:6656];
        1241: state_byte <= hashes[6655:6648];
        1242: state_byte <= hashes[6647:6640];
        1243: state_byte <= hashes[6639:6632];
        1244: state_byte <= hashes[6631:6624];
        1245: state_byte <= hashes[6623:6616];
        1246: state_byte <= hashes[6615:6608];
        1247: state_byte <= hashes[6607:6600];
        1248: state_byte <= hashes[6599:6592];
        1249: state_byte <= hashes[6591:6584];
        1250: state_byte <= hashes[6583:6576];
        1251: state_byte <= hashes[6575:6568];
        1252: state_byte <= hashes[6567:6560];
        1253: state_byte <= hashes[6559:6552];
        1254: state_byte <= hashes[6551:6544];
        1255: state_byte <= hashes[6543:6536];
        1256: state_byte <= hashes[6535:6528];
        1257: state_byte <= hashes[6527:6520];
        1258: state_byte <= hashes[6519:6512];
        1259: state_byte <= hashes[6511:6504];
        1260: state_byte <= hashes[6503:6496];
        1261: state_byte <= hashes[6495:6488];
        1262: state_byte <= hashes[6487:6480];
        1263: state_byte <= hashes[6479:6472];
        1264: state_byte <= hashes[6471:6464];
        1265: state_byte <= hashes[6463:6456];
        1266: state_byte <= hashes[6455:6448];
        1267: state_byte <= hashes[6447:6440];
        1268: state_byte <= hashes[6439:6432];
        1269: state_byte <= hashes[6431:6424];
        1270: state_byte <= hashes[6423:6416];
        1271: state_byte <= hashes[6415:6408];
        1272: state_byte <= hashes[6407:6400];
        1273: state_byte <= hashes[6399:6392];
        1274: state_byte <= hashes[6391:6384];
        1275: state_byte <= hashes[6383:6376];
        1276: state_byte <= hashes[6375:6368];
        1277: state_byte <= hashes[6367:6360];
        1278: state_byte <= hashes[6359:6352];
        1279: state_byte <= hashes[6351:6344];
        1280: state_byte <= hashes[6343:6336];
        1281: state_byte <= hashes[6335:6328];
        1282: state_byte <= hashes[6327:6320];
        1283: state_byte <= hashes[6319:6312];
        1284: state_byte <= hashes[6311:6304];
        1285: state_byte <= hashes[6303:6296];
        1286: state_byte <= hashes[6295:6288];
        1287: state_byte <= hashes[6287:6280];
        1288: state_byte <= hashes[6279:6272];
        1289: state_byte <= hashes[6271:6264];
        1290: state_byte <= hashes[6263:6256];
        1291: state_byte <= hashes[6255:6248];
        1292: state_byte <= hashes[6247:6240];
        1293: state_byte <= hashes[6239:6232];
        1294: state_byte <= hashes[6231:6224];
        1295: state_byte <= hashes[6223:6216];
        1296: state_byte <= hashes[6215:6208];
        1297: state_byte <= hashes[6207:6200];
        1298: state_byte <= hashes[6199:6192];
        1299: state_byte <= hashes[6191:6184];
        1300: state_byte <= hashes[6183:6176];
        1301: state_byte <= hashes[6175:6168];
        1302: state_byte <= hashes[6167:6160];
        1303: state_byte <= hashes[6159:6152];
        1304: state_byte <= hashes[6151:6144];
        1305: state_byte <= hashes[6143:6136];
        1306: state_byte <= hashes[6135:6128];
        1307: state_byte <= hashes[6127:6120];
        1308: state_byte <= hashes[6119:6112];
        1309: state_byte <= hashes[6111:6104];
        1310: state_byte <= hashes[6103:6096];
        1311: state_byte <= hashes[6095:6088];
        1312: state_byte <= hashes[6087:6080];
        1313: state_byte <= hashes[6079:6072];
        1314: state_byte <= hashes[6071:6064];
        1315: state_byte <= hashes[6063:6056];
        1316: state_byte <= hashes[6055:6048];
        1317: state_byte <= hashes[6047:6040];
        1318: state_byte <= hashes[6039:6032];
        1319: state_byte <= hashes[6031:6024];
        1320: state_byte <= hashes[6023:6016];
        1321: state_byte <= hashes[6015:6008];
        1322: state_byte <= hashes[6007:6000];
        1323: state_byte <= hashes[5999:5992];
        1324: state_byte <= hashes[5991:5984];
        1325: state_byte <= hashes[5983:5976];
        1326: state_byte <= hashes[5975:5968];
        1327: state_byte <= hashes[5967:5960];
        1328: state_byte <= hashes[5959:5952];
        1329: state_byte <= hashes[5951:5944];
        1330: state_byte <= hashes[5943:5936];
        1331: state_byte <= hashes[5935:5928];
        1332: state_byte <= hashes[5927:5920];
        1333: state_byte <= hashes[5919:5912];
        1334: state_byte <= hashes[5911:5904];
        1335: state_byte <= hashes[5903:5896];
        1336: state_byte <= hashes[5895:5888];
        1337: state_byte <= hashes[5887:5880];
        1338: state_byte <= hashes[5879:5872];
        1339: state_byte <= hashes[5871:5864];
        1340: state_byte <= hashes[5863:5856];
        1341: state_byte <= hashes[5855:5848];
        1342: state_byte <= hashes[5847:5840];
        1343: state_byte <= hashes[5839:5832];
        1344: state_byte <= hashes[5831:5824];
        1345: state_byte <= hashes[5823:5816];
        1346: state_byte <= hashes[5815:5808];
        1347: state_byte <= hashes[5807:5800];
        1348: state_byte <= hashes[5799:5792];
        1349: state_byte <= hashes[5791:5784];
        1350: state_byte <= hashes[5783:5776];
        1351: state_byte <= hashes[5775:5768];
        1352: state_byte <= hashes[5767:5760];
        1353: state_byte <= hashes[5759:5752];
        1354: state_byte <= hashes[5751:5744];
        1355: state_byte <= hashes[5743:5736];
        1356: state_byte <= hashes[5735:5728];
        1357: state_byte <= hashes[5727:5720];
        1358: state_byte <= hashes[5719:5712];
        1359: state_byte <= hashes[5711:5704];
        1360: state_byte <= hashes[5703:5696];
        1361: state_byte <= hashes[5695:5688];
        1362: state_byte <= hashes[5687:5680];
        1363: state_byte <= hashes[5679:5672];
        1364: state_byte <= hashes[5671:5664];
        1365: state_byte <= hashes[5663:5656];
        1366: state_byte <= hashes[5655:5648];
        1367: state_byte <= hashes[5647:5640];
        1368: state_byte <= hashes[5639:5632];
        1369: state_byte <= hashes[5631:5624];
        1370: state_byte <= hashes[5623:5616];
        1371: state_byte <= hashes[5615:5608];
        1372: state_byte <= hashes[5607:5600];
        1373: state_byte <= hashes[5599:5592];
        1374: state_byte <= hashes[5591:5584];
        1375: state_byte <= hashes[5583:5576];
        1376: state_byte <= hashes[5575:5568];
        1377: state_byte <= hashes[5567:5560];
        1378: state_byte <= hashes[5559:5552];
        1379: state_byte <= hashes[5551:5544];
        1380: state_byte <= hashes[5543:5536];
        1381: state_byte <= hashes[5535:5528];
        1382: state_byte <= hashes[5527:5520];
        1383: state_byte <= hashes[5519:5512];
        1384: state_byte <= hashes[5511:5504];
        1385: state_byte <= hashes[5503:5496];
        1386: state_byte <= hashes[5495:5488];
        1387: state_byte <= hashes[5487:5480];
        1388: state_byte <= hashes[5479:5472];
        1389: state_byte <= hashes[5471:5464];
        1390: state_byte <= hashes[5463:5456];
        1391: state_byte <= hashes[5455:5448];
        1392: state_byte <= hashes[5447:5440];
        1393: state_byte <= hashes[5439:5432];
        1394: state_byte <= hashes[5431:5424];
        1395: state_byte <= hashes[5423:5416];
        1396: state_byte <= hashes[5415:5408];
        1397: state_byte <= hashes[5407:5400];
        1398: state_byte <= hashes[5399:5392];
        1399: state_byte <= hashes[5391:5384];
        1400: state_byte <= hashes[5383:5376];
        1401: state_byte <= hashes[5375:5368];
        1402: state_byte <= hashes[5367:5360];
        1403: state_byte <= hashes[5359:5352];
        1404: state_byte <= hashes[5351:5344];
        1405: state_byte <= hashes[5343:5336];
        1406: state_byte <= hashes[5335:5328];
        1407: state_byte <= hashes[5327:5320];
        1408: state_byte <= hashes[5319:5312];
        1409: state_byte <= hashes[5311:5304];
        1410: state_byte <= hashes[5303:5296];
        1411: state_byte <= hashes[5295:5288];
        1412: state_byte <= hashes[5287:5280];
        1413: state_byte <= hashes[5279:5272];
        1414: state_byte <= hashes[5271:5264];
        1415: state_byte <= hashes[5263:5256];
        1416: state_byte <= hashes[5255:5248];
        1417: state_byte <= hashes[5247:5240];
        1418: state_byte <= hashes[5239:5232];
        1419: state_byte <= hashes[5231:5224];
        1420: state_byte <= hashes[5223:5216];
        1421: state_byte <= hashes[5215:5208];
        1422: state_byte <= hashes[5207:5200];
        1423: state_byte <= hashes[5199:5192];
        1424: state_byte <= hashes[5191:5184];
        1425: state_byte <= hashes[5183:5176];
        1426: state_byte <= hashes[5175:5168];
        1427: state_byte <= hashes[5167:5160];
        1428: state_byte <= hashes[5159:5152];
        1429: state_byte <= hashes[5151:5144];
        1430: state_byte <= hashes[5143:5136];
        1431: state_byte <= hashes[5135:5128];
        1432: state_byte <= hashes[5127:5120];
        1433: state_byte <= hashes[5119:5112];
        1434: state_byte <= hashes[5111:5104];
        1435: state_byte <= hashes[5103:5096];
        1436: state_byte <= hashes[5095:5088];
        1437: state_byte <= hashes[5087:5080];
        1438: state_byte <= hashes[5079:5072];
        1439: state_byte <= hashes[5071:5064];
        1440: state_byte <= hashes[5063:5056];
        1441: state_byte <= hashes[5055:5048];
        1442: state_byte <= hashes[5047:5040];
        1443: state_byte <= hashes[5039:5032];
        1444: state_byte <= hashes[5031:5024];
        1445: state_byte <= hashes[5023:5016];
        1446: state_byte <= hashes[5015:5008];
        1447: state_byte <= hashes[5007:5000];
        1448: state_byte <= hashes[4999:4992];
        1449: state_byte <= hashes[4991:4984];
        1450: state_byte <= hashes[4983:4976];
        1451: state_byte <= hashes[4975:4968];
        1452: state_byte <= hashes[4967:4960];
        1453: state_byte <= hashes[4959:4952];
        1454: state_byte <= hashes[4951:4944];
        1455: state_byte <= hashes[4943:4936];
        1456: state_byte <= hashes[4935:4928];
        1457: state_byte <= hashes[4927:4920];
        1458: state_byte <= hashes[4919:4912];
        1459: state_byte <= hashes[4911:4904];
        1460: state_byte <= hashes[4903:4896];
        1461: state_byte <= hashes[4895:4888];
        1462: state_byte <= hashes[4887:4880];
        1463: state_byte <= hashes[4879:4872];
        1464: state_byte <= hashes[4871:4864];
        1465: state_byte <= hashes[4863:4856];
        1466: state_byte <= hashes[4855:4848];
        1467: state_byte <= hashes[4847:4840];
        1468: state_byte <= hashes[4839:4832];
        1469: state_byte <= hashes[4831:4824];
        1470: state_byte <= hashes[4823:4816];
        1471: state_byte <= hashes[4815:4808];
        1472: state_byte <= hashes[4807:4800];
        1473: state_byte <= hashes[4799:4792];
        1474: state_byte <= hashes[4791:4784];
        1475: state_byte <= hashes[4783:4776];
        1476: state_byte <= hashes[4775:4768];
        1477: state_byte <= hashes[4767:4760];
        1478: state_byte <= hashes[4759:4752];
        1479: state_byte <= hashes[4751:4744];
        1480: state_byte <= hashes[4743:4736];
        1481: state_byte <= hashes[4735:4728];
        1482: state_byte <= hashes[4727:4720];
        1483: state_byte <= hashes[4719:4712];
        1484: state_byte <= hashes[4711:4704];
        1485: state_byte <= hashes[4703:4696];
        1486: state_byte <= hashes[4695:4688];
        1487: state_byte <= hashes[4687:4680];
        1488: state_byte <= hashes[4679:4672];
        1489: state_byte <= hashes[4671:4664];
        1490: state_byte <= hashes[4663:4656];
        1491: state_byte <= hashes[4655:4648];
        1492: state_byte <= hashes[4647:4640];
        1493: state_byte <= hashes[4639:4632];
        1494: state_byte <= hashes[4631:4624];
        1495: state_byte <= hashes[4623:4616];
        1496: state_byte <= hashes[4615:4608];
        1497: state_byte <= hashes[4607:4600];
        1498: state_byte <= hashes[4599:4592];
        1499: state_byte <= hashes[4591:4584];
        1500: state_byte <= hashes[4583:4576];
        1501: state_byte <= hashes[4575:4568];
        1502: state_byte <= hashes[4567:4560];
        1503: state_byte <= hashes[4559:4552];
        1504: state_byte <= hashes[4551:4544];
        1505: state_byte <= hashes[4543:4536];
        1506: state_byte <= hashes[4535:4528];
        1507: state_byte <= hashes[4527:4520];
        1508: state_byte <= hashes[4519:4512];
        1509: state_byte <= hashes[4511:4504];
        1510: state_byte <= hashes[4503:4496];
        1511: state_byte <= hashes[4495:4488];
        1512: state_byte <= hashes[4487:4480];
        1513: state_byte <= hashes[4479:4472];
        1514: state_byte <= hashes[4471:4464];
        1515: state_byte <= hashes[4463:4456];
        1516: state_byte <= hashes[4455:4448];
        1517: state_byte <= hashes[4447:4440];
        1518: state_byte <= hashes[4439:4432];
        1519: state_byte <= hashes[4431:4424];
        1520: state_byte <= hashes[4423:4416];
        1521: state_byte <= hashes[4415:4408];
        1522: state_byte <= hashes[4407:4400];
        1523: state_byte <= hashes[4399:4392];
        1524: state_byte <= hashes[4391:4384];
        1525: state_byte <= hashes[4383:4376];
        1526: state_byte <= hashes[4375:4368];
        1527: state_byte <= hashes[4367:4360];
        1528: state_byte <= hashes[4359:4352];
        1529: state_byte <= hashes[4351:4344];
        1530: state_byte <= hashes[4343:4336];
        1531: state_byte <= hashes[4335:4328];
        1532: state_byte <= hashes[4327:4320];
        1533: state_byte <= hashes[4319:4312];
        1534: state_byte <= hashes[4311:4304];
        1535: state_byte <= hashes[4303:4296];
        1536: state_byte <= hashes[4295:4288];
        1537: state_byte <= hashes[4287:4280];
        1538: state_byte <= hashes[4279:4272];
        1539: state_byte <= hashes[4271:4264];
        1540: state_byte <= hashes[4263:4256];
        1541: state_byte <= hashes[4255:4248];
        1542: state_byte <= hashes[4247:4240];
        1543: state_byte <= hashes[4239:4232];
        1544: state_byte <= hashes[4231:4224];
        1545: state_byte <= hashes[4223:4216];
        1546: state_byte <= hashes[4215:4208];
        1547: state_byte <= hashes[4207:4200];
        1548: state_byte <= hashes[4199:4192];
        1549: state_byte <= hashes[4191:4184];
        1550: state_byte <= hashes[4183:4176];
        1551: state_byte <= hashes[4175:4168];
        1552: state_byte <= hashes[4167:4160];
        1553: state_byte <= hashes[4159:4152];
        1554: state_byte <= hashes[4151:4144];
        1555: state_byte <= hashes[4143:4136];
        1556: state_byte <= hashes[4135:4128];
        1557: state_byte <= hashes[4127:4120];
        1558: state_byte <= hashes[4119:4112];
        1559: state_byte <= hashes[4111:4104];
        1560: state_byte <= hashes[4103:4096];
        1561: state_byte <= hashes[4095:4088];
        1562: state_byte <= hashes[4087:4080];
        1563: state_byte <= hashes[4079:4072];
        1564: state_byte <= hashes[4071:4064];
        1565: state_byte <= hashes[4063:4056];
        1566: state_byte <= hashes[4055:4048];
        1567: state_byte <= hashes[4047:4040];
        1568: state_byte <= hashes[4039:4032];
        1569: state_byte <= hashes[4031:4024];
        1570: state_byte <= hashes[4023:4016];
        1571: state_byte <= hashes[4015:4008];
        1572: state_byte <= hashes[4007:4000];
        1573: state_byte <= hashes[3999:3992];
        1574: state_byte <= hashes[3991:3984];
        1575: state_byte <= hashes[3983:3976];
        1576: state_byte <= hashes[3975:3968];
        1577: state_byte <= hashes[3967:3960];
        1578: state_byte <= hashes[3959:3952];
        1579: state_byte <= hashes[3951:3944];
        1580: state_byte <= hashes[3943:3936];
        1581: state_byte <= hashes[3935:3928];
        1582: state_byte <= hashes[3927:3920];
        1583: state_byte <= hashes[3919:3912];
        1584: state_byte <= hashes[3911:3904];
        1585: state_byte <= hashes[3903:3896];
        1586: state_byte <= hashes[3895:3888];
        1587: state_byte <= hashes[3887:3880];
        1588: state_byte <= hashes[3879:3872];
        1589: state_byte <= hashes[3871:3864];
        1590: state_byte <= hashes[3863:3856];
        1591: state_byte <= hashes[3855:3848];
        1592: state_byte <= hashes[3847:3840];
        1593: state_byte <= hashes[3839:3832];
        1594: state_byte <= hashes[3831:3824];
        1595: state_byte <= hashes[3823:3816];
        1596: state_byte <= hashes[3815:3808];
        1597: state_byte <= hashes[3807:3800];
        1598: state_byte <= hashes[3799:3792];
        1599: state_byte <= hashes[3791:3784];
        1600: state_byte <= hashes[3783:3776];
        1601: state_byte <= hashes[3775:3768];
        1602: state_byte <= hashes[3767:3760];
        1603: state_byte <= hashes[3759:3752];
        1604: state_byte <= hashes[3751:3744];
        1605: state_byte <= hashes[3743:3736];
        1606: state_byte <= hashes[3735:3728];
        1607: state_byte <= hashes[3727:3720];
        1608: state_byte <= hashes[3719:3712];
        1609: state_byte <= hashes[3711:3704];
        1610: state_byte <= hashes[3703:3696];
        1611: state_byte <= hashes[3695:3688];
        1612: state_byte <= hashes[3687:3680];
        1613: state_byte <= hashes[3679:3672];
        1614: state_byte <= hashes[3671:3664];
        1615: state_byte <= hashes[3663:3656];
        1616: state_byte <= hashes[3655:3648];
        1617: state_byte <= hashes[3647:3640];
        1618: state_byte <= hashes[3639:3632];
        1619: state_byte <= hashes[3631:3624];
        1620: state_byte <= hashes[3623:3616];
        1621: state_byte <= hashes[3615:3608];
        1622: state_byte <= hashes[3607:3600];
        1623: state_byte <= hashes[3599:3592];
        1624: state_byte <= hashes[3591:3584];
        1625: state_byte <= hashes[3583:3576];
        1626: state_byte <= hashes[3575:3568];
        1627: state_byte <= hashes[3567:3560];
        1628: state_byte <= hashes[3559:3552];
        1629: state_byte <= hashes[3551:3544];
        1630: state_byte <= hashes[3543:3536];
        1631: state_byte <= hashes[3535:3528];
        1632: state_byte <= hashes[3527:3520];
        1633: state_byte <= hashes[3519:3512];
        1634: state_byte <= hashes[3511:3504];
        1635: state_byte <= hashes[3503:3496];
        1636: state_byte <= hashes[3495:3488];
        1637: state_byte <= hashes[3487:3480];
        1638: state_byte <= hashes[3479:3472];
        1639: state_byte <= hashes[3471:3464];
        1640: state_byte <= hashes[3463:3456];
        1641: state_byte <= hashes[3455:3448];
        1642: state_byte <= hashes[3447:3440];
        1643: state_byte <= hashes[3439:3432];
        1644: state_byte <= hashes[3431:3424];
        1645: state_byte <= hashes[3423:3416];
        1646: state_byte <= hashes[3415:3408];
        1647: state_byte <= hashes[3407:3400];
        1648: state_byte <= hashes[3399:3392];
        1649: state_byte <= hashes[3391:3384];
        1650: state_byte <= hashes[3383:3376];
        1651: state_byte <= hashes[3375:3368];
        1652: state_byte <= hashes[3367:3360];
        1653: state_byte <= hashes[3359:3352];
        1654: state_byte <= hashes[3351:3344];
        1655: state_byte <= hashes[3343:3336];
        1656: state_byte <= hashes[3335:3328];
        1657: state_byte <= hashes[3327:3320];
        1658: state_byte <= hashes[3319:3312];
        1659: state_byte <= hashes[3311:3304];
        1660: state_byte <= hashes[3303:3296];
        1661: state_byte <= hashes[3295:3288];
        1662: state_byte <= hashes[3287:3280];
        1663: state_byte <= hashes[3279:3272];
        1664: state_byte <= hashes[3271:3264];
        1665: state_byte <= hashes[3263:3256];
        1666: state_byte <= hashes[3255:3248];
        1667: state_byte <= hashes[3247:3240];
        1668: state_byte <= hashes[3239:3232];
        1669: state_byte <= hashes[3231:3224];
        1670: state_byte <= hashes[3223:3216];
        1671: state_byte <= hashes[3215:3208];
        1672: state_byte <= hashes[3207:3200];
        1673: state_byte <= hashes[3199:3192];
        1674: state_byte <= hashes[3191:3184];
        1675: state_byte <= hashes[3183:3176];
        1676: state_byte <= hashes[3175:3168];
        1677: state_byte <= hashes[3167:3160];
        1678: state_byte <= hashes[3159:3152];
        1679: state_byte <= hashes[3151:3144];
        1680: state_byte <= hashes[3143:3136];
        1681: state_byte <= hashes[3135:3128];
        1682: state_byte <= hashes[3127:3120];
        1683: state_byte <= hashes[3119:3112];
        1684: state_byte <= hashes[3111:3104];
        1685: state_byte <= hashes[3103:3096];
        1686: state_byte <= hashes[3095:3088];
        1687: state_byte <= hashes[3087:3080];
        1688: state_byte <= hashes[3079:3072];
        1689: state_byte <= hashes[3071:3064];
        1690: state_byte <= hashes[3063:3056];
        1691: state_byte <= hashes[3055:3048];
        1692: state_byte <= hashes[3047:3040];
        1693: state_byte <= hashes[3039:3032];
        1694: state_byte <= hashes[3031:3024];
        1695: state_byte <= hashes[3023:3016];
        1696: state_byte <= hashes[3015:3008];
        1697: state_byte <= hashes[3007:3000];
        1698: state_byte <= hashes[2999:2992];
        1699: state_byte <= hashes[2991:2984];
        1700: state_byte <= hashes[2983:2976];
        1701: state_byte <= hashes[2975:2968];
        1702: state_byte <= hashes[2967:2960];
        1703: state_byte <= hashes[2959:2952];
        1704: state_byte <= hashes[2951:2944];
        1705: state_byte <= hashes[2943:2936];
        1706: state_byte <= hashes[2935:2928];
        1707: state_byte <= hashes[2927:2920];
        1708: state_byte <= hashes[2919:2912];
        1709: state_byte <= hashes[2911:2904];
        1710: state_byte <= hashes[2903:2896];
        1711: state_byte <= hashes[2895:2888];
        1712: state_byte <= hashes[2887:2880];
        1713: state_byte <= hashes[2879:2872];
        1714: state_byte <= hashes[2871:2864];
        1715: state_byte <= hashes[2863:2856];
        1716: state_byte <= hashes[2855:2848];
        1717: state_byte <= hashes[2847:2840];
        1718: state_byte <= hashes[2839:2832];
        1719: state_byte <= hashes[2831:2824];
        1720: state_byte <= hashes[2823:2816];
        1721: state_byte <= hashes[2815:2808];
        1722: state_byte <= hashes[2807:2800];
        1723: state_byte <= hashes[2799:2792];
        1724: state_byte <= hashes[2791:2784];
        1725: state_byte <= hashes[2783:2776];
        1726: state_byte <= hashes[2775:2768];
        1727: state_byte <= hashes[2767:2760];
        1728: state_byte <= hashes[2759:2752];
        1729: state_byte <= hashes[2751:2744];
        1730: state_byte <= hashes[2743:2736];
        1731: state_byte <= hashes[2735:2728];
        1732: state_byte <= hashes[2727:2720];
        1733: state_byte <= hashes[2719:2712];
        1734: state_byte <= hashes[2711:2704];
        1735: state_byte <= hashes[2703:2696];
        1736: state_byte <= hashes[2695:2688];
        1737: state_byte <= hashes[2687:2680];
        1738: state_byte <= hashes[2679:2672];
        1739: state_byte <= hashes[2671:2664];
        1740: state_byte <= hashes[2663:2656];
        1741: state_byte <= hashes[2655:2648];
        1742: state_byte <= hashes[2647:2640];
        1743: state_byte <= hashes[2639:2632];
        1744: state_byte <= hashes[2631:2624];
        1745: state_byte <= hashes[2623:2616];
        1746: state_byte <= hashes[2615:2608];
        1747: state_byte <= hashes[2607:2600];
        1748: state_byte <= hashes[2599:2592];
        1749: state_byte <= hashes[2591:2584];
        1750: state_byte <= hashes[2583:2576];
        1751: state_byte <= hashes[2575:2568];
        1752: state_byte <= hashes[2567:2560];
        1753: state_byte <= hashes[2559:2552];
        1754: state_byte <= hashes[2551:2544];
        1755: state_byte <= hashes[2543:2536];
        1756: state_byte <= hashes[2535:2528];
        1757: state_byte <= hashes[2527:2520];
        1758: state_byte <= hashes[2519:2512];
        1759: state_byte <= hashes[2511:2504];
        1760: state_byte <= hashes[2503:2496];
        1761: state_byte <= hashes[2495:2488];
        1762: state_byte <= hashes[2487:2480];
        1763: state_byte <= hashes[2479:2472];
        1764: state_byte <= hashes[2471:2464];
        1765: state_byte <= hashes[2463:2456];
        1766: state_byte <= hashes[2455:2448];
        1767: state_byte <= hashes[2447:2440];
        1768: state_byte <= hashes[2439:2432];
        1769: state_byte <= hashes[2431:2424];
        1770: state_byte <= hashes[2423:2416];
        1771: state_byte <= hashes[2415:2408];
        1772: state_byte <= hashes[2407:2400];
        1773: state_byte <= hashes[2399:2392];
        1774: state_byte <= hashes[2391:2384];
        1775: state_byte <= hashes[2383:2376];
        1776: state_byte <= hashes[2375:2368];
        1777: state_byte <= hashes[2367:2360];
        1778: state_byte <= hashes[2359:2352];
        1779: state_byte <= hashes[2351:2344];
        1780: state_byte <= hashes[2343:2336];
        1781: state_byte <= hashes[2335:2328];
        1782: state_byte <= hashes[2327:2320];
        1783: state_byte <= hashes[2319:2312];
        1784: state_byte <= hashes[2311:2304];
        1785: state_byte <= hashes[2303:2296];
        1786: state_byte <= hashes[2295:2288];
        1787: state_byte <= hashes[2287:2280];
        1788: state_byte <= hashes[2279:2272];
        1789: state_byte <= hashes[2271:2264];
        1790: state_byte <= hashes[2263:2256];
        1791: state_byte <= hashes[2255:2248];
        1792: state_byte <= hashes[2247:2240];
        1793: state_byte <= hashes[2239:2232];
        1794: state_byte <= hashes[2231:2224];
        1795: state_byte <= hashes[2223:2216];
        1796: state_byte <= hashes[2215:2208];
        1797: state_byte <= hashes[2207:2200];
        1798: state_byte <= hashes[2199:2192];
        1799: state_byte <= hashes[2191:2184];
        1800: state_byte <= hashes[2183:2176];
        1801: state_byte <= hashes[2175:2168];
        1802: state_byte <= hashes[2167:2160];
        1803: state_byte <= hashes[2159:2152];
        1804: state_byte <= hashes[2151:2144];
        1805: state_byte <= hashes[2143:2136];
        1806: state_byte <= hashes[2135:2128];
        1807: state_byte <= hashes[2127:2120];
        1808: state_byte <= hashes[2119:2112];
        1809: state_byte <= hashes[2111:2104];
        1810: state_byte <= hashes[2103:2096];
        1811: state_byte <= hashes[2095:2088];
        1812: state_byte <= hashes[2087:2080];
        1813: state_byte <= hashes[2079:2072];
        1814: state_byte <= hashes[2071:2064];
        1815: state_byte <= hashes[2063:2056];
        1816: state_byte <= hashes[2055:2048];
        1817: state_byte <= hashes[2047:2040];
        1818: state_byte <= hashes[2039:2032];
        1819: state_byte <= hashes[2031:2024];
        1820: state_byte <= hashes[2023:2016];
        1821: state_byte <= hashes[2015:2008];
        1822: state_byte <= hashes[2007:2000];
        1823: state_byte <= hashes[1999:1992];
        1824: state_byte <= hashes[1991:1984];
        1825: state_byte <= hashes[1983:1976];
        1826: state_byte <= hashes[1975:1968];
        1827: state_byte <= hashes[1967:1960];
        1828: state_byte <= hashes[1959:1952];
        1829: state_byte <= hashes[1951:1944];
        1830: state_byte <= hashes[1943:1936];
        1831: state_byte <= hashes[1935:1928];
        1832: state_byte <= hashes[1927:1920];
        1833: state_byte <= hashes[1919:1912];
        1834: state_byte <= hashes[1911:1904];
        1835: state_byte <= hashes[1903:1896];
        1836: state_byte <= hashes[1895:1888];
        1837: state_byte <= hashes[1887:1880];
        1838: state_byte <= hashes[1879:1872];
        1839: state_byte <= hashes[1871:1864];
        1840: state_byte <= hashes[1863:1856];
        1841: state_byte <= hashes[1855:1848];
        1842: state_byte <= hashes[1847:1840];
        1843: state_byte <= hashes[1839:1832];
        1844: state_byte <= hashes[1831:1824];
        1845: state_byte <= hashes[1823:1816];
        1846: state_byte <= hashes[1815:1808];
        1847: state_byte <= hashes[1807:1800];
        1848: state_byte <= hashes[1799:1792];
        1849: state_byte <= hashes[1791:1784];
        1850: state_byte <= hashes[1783:1776];
        1851: state_byte <= hashes[1775:1768];
        1852: state_byte <= hashes[1767:1760];
        1853: state_byte <= hashes[1759:1752];
        1854: state_byte <= hashes[1751:1744];
        1855: state_byte <= hashes[1743:1736];
        1856: state_byte <= hashes[1735:1728];
        1857: state_byte <= hashes[1727:1720];
        1858: state_byte <= hashes[1719:1712];
        1859: state_byte <= hashes[1711:1704];
        1860: state_byte <= hashes[1703:1696];
        1861: state_byte <= hashes[1695:1688];
        1862: state_byte <= hashes[1687:1680];
        1863: state_byte <= hashes[1679:1672];
        1864: state_byte <= hashes[1671:1664];
        1865: state_byte <= hashes[1663:1656];
        1866: state_byte <= hashes[1655:1648];
        1867: state_byte <= hashes[1647:1640];
        1868: state_byte <= hashes[1639:1632];
        1869: state_byte <= hashes[1631:1624];
        1870: state_byte <= hashes[1623:1616];
        1871: state_byte <= hashes[1615:1608];
        1872: state_byte <= hashes[1607:1600];
        1873: state_byte <= hashes[1599:1592];
        1874: state_byte <= hashes[1591:1584];
        1875: state_byte <= hashes[1583:1576];
        1876: state_byte <= hashes[1575:1568];
        1877: state_byte <= hashes[1567:1560];
        1878: state_byte <= hashes[1559:1552];
        1879: state_byte <= hashes[1551:1544];
        1880: state_byte <= hashes[1543:1536];
        1881: state_byte <= hashes[1535:1528];
        1882: state_byte <= hashes[1527:1520];
        1883: state_byte <= hashes[1519:1512];
        1884: state_byte <= hashes[1511:1504];
        1885: state_byte <= hashes[1503:1496];
        1886: state_byte <= hashes[1495:1488];
        1887: state_byte <= hashes[1487:1480];
        1888: state_byte <= hashes[1479:1472];
        1889: state_byte <= hashes[1471:1464];
        1890: state_byte <= hashes[1463:1456];
        1891: state_byte <= hashes[1455:1448];
        1892: state_byte <= hashes[1447:1440];
        1893: state_byte <= hashes[1439:1432];
        1894: state_byte <= hashes[1431:1424];
        1895: state_byte <= hashes[1423:1416];
        1896: state_byte <= hashes[1415:1408];
        1897: state_byte <= hashes[1407:1400];
        1898: state_byte <= hashes[1399:1392];
        1899: state_byte <= hashes[1391:1384];
        1900: state_byte <= hashes[1383:1376];
        1901: state_byte <= hashes[1375:1368];
        1902: state_byte <= hashes[1367:1360];
        1903: state_byte <= hashes[1359:1352];
        1904: state_byte <= hashes[1351:1344];
        1905: state_byte <= hashes[1343:1336];
        1906: state_byte <= hashes[1335:1328];
        1907: state_byte <= hashes[1327:1320];
        1908: state_byte <= hashes[1319:1312];
        1909: state_byte <= hashes[1311:1304];
        1910: state_byte <= hashes[1303:1296];
        1911: state_byte <= hashes[1295:1288];
        1912: state_byte <= hashes[1287:1280];
        1913: state_byte <= hashes[1279:1272];
        1914: state_byte <= hashes[1271:1264];
        1915: state_byte <= hashes[1263:1256];
        1916: state_byte <= hashes[1255:1248];
        1917: state_byte <= hashes[1247:1240];
        1918: state_byte <= hashes[1239:1232];
        1919: state_byte <= hashes[1231:1224];
        1920: state_byte <= hashes[1223:1216];
        1921: state_byte <= hashes[1215:1208];
        1922: state_byte <= hashes[1207:1200];
        1923: state_byte <= hashes[1199:1192];
        1924: state_byte <= hashes[1191:1184];
        1925: state_byte <= hashes[1183:1176];
        1926: state_byte <= hashes[1175:1168];
        1927: state_byte <= hashes[1167:1160];
        1928: state_byte <= hashes[1159:1152];
        1929: state_byte <= hashes[1151:1144];
        1930: state_byte <= hashes[1143:1136];
        1931: state_byte <= hashes[1135:1128];
        1932: state_byte <= hashes[1127:1120];
        1933: state_byte <= hashes[1119:1112];
        1934: state_byte <= hashes[1111:1104];
        1935: state_byte <= hashes[1103:1096];
        1936: state_byte <= hashes[1095:1088];
        1937: state_byte <= hashes[1087:1080];
        1938: state_byte <= hashes[1079:1072];
        1939: state_byte <= hashes[1071:1064];
        1940: state_byte <= hashes[1063:1056];
        1941: state_byte <= hashes[1055:1048];
        1942: state_byte <= hashes[1047:1040];
        1943: state_byte <= hashes[1039:1032];
        1944: state_byte <= hashes[1031:1024];
        1945: state_byte <= hashes[1023:1016];
        1946: state_byte <= hashes[1015:1008];
        1947: state_byte <= hashes[1007:1000];
        1948: state_byte <= hashes[999:992];
        1949: state_byte <= hashes[991:984];
        1950: state_byte <= hashes[983:976];
        1951: state_byte <= hashes[975:968];
        1952: state_byte <= hashes[967:960];
        1953: state_byte <= hashes[959:952];
        1954: state_byte <= hashes[951:944];
        1955: state_byte <= hashes[943:936];
        1956: state_byte <= hashes[935:928];
        1957: state_byte <= hashes[927:920];
        1958: state_byte <= hashes[919:912];
        1959: state_byte <= hashes[911:904];
        1960: state_byte <= hashes[903:896];
        1961: state_byte <= hashes[895:888];
        1962: state_byte <= hashes[887:880];
        1963: state_byte <= hashes[879:872];
        1964: state_byte <= hashes[871:864];
        1965: state_byte <= hashes[863:856];
        1966: state_byte <= hashes[855:848];
        1967: state_byte <= hashes[847:840];
        1968: state_byte <= hashes[839:832];
        1969: state_byte <= hashes[831:824];
        1970: state_byte <= hashes[823:816];
        1971: state_byte <= hashes[815:808];
        1972: state_byte <= hashes[807:800];
        1973: state_byte <= hashes[799:792];
        1974: state_byte <= hashes[791:784];
        1975: state_byte <= hashes[783:776];
        1976: state_byte <= hashes[775:768];
        1977: state_byte <= hashes[767:760];
        1978: state_byte <= hashes[759:752];
        1979: state_byte <= hashes[751:744];
        1980: state_byte <= hashes[743:736];
        1981: state_byte <= hashes[735:728];
        1982: state_byte <= hashes[727:720];
        1983: state_byte <= hashes[719:712];
        1984: state_byte <= hashes[711:704];
        1985: state_byte <= hashes[703:696];
        1986: state_byte <= hashes[695:688];
        1987: state_byte <= hashes[687:680];
        1988: state_byte <= hashes[679:672];
        1989: state_byte <= hashes[671:664];
        1990: state_byte <= hashes[663:656];
        1991: state_byte <= hashes[655:648];
        1992: state_byte <= hashes[647:640];
        1993: state_byte <= hashes[639:632];
        1994: state_byte <= hashes[631:624];
        1995: state_byte <= hashes[623:616];
        1996: state_byte <= hashes[615:608];
        1997: state_byte <= hashes[607:600];
        1998: state_byte <= hashes[599:592];
        1999: state_byte <= hashes[591:584];
        2000: state_byte <= hashes[583:576];
        2001: state_byte <= hashes[575:568];
        2002: state_byte <= hashes[567:560];
        2003: state_byte <= hashes[559:552];
        2004: state_byte <= hashes[551:544];
        2005: state_byte <= hashes[543:536];
        2006: state_byte <= hashes[535:528];
        2007: state_byte <= hashes[527:520];
        2008: state_byte <= hashes[519:512];
        2009: state_byte <= hashes[511:504];
        2010: state_byte <= hashes[503:496];
        2011: state_byte <= hashes[495:488];
        2012: state_byte <= hashes[487:480];
        2013: state_byte <= hashes[479:472];
        2014: state_byte <= hashes[471:464];
        2015: state_byte <= hashes[463:456];
        2016: state_byte <= hashes[455:448];
        2017: state_byte <= hashes[447:440];
        2018: state_byte <= hashes[439:432];
        2019: state_byte <= hashes[431:424];
        2020: state_byte <= hashes[423:416];
        2021: state_byte <= hashes[415:408];
        2022: state_byte <= hashes[407:400];
        2023: state_byte <= hashes[399:392];
        2024: state_byte <= hashes[391:384];
        2025: state_byte <= hashes[383:376];
        2026: state_byte <= hashes[375:368];
        2027: state_byte <= hashes[367:360];
        2028: state_byte <= hashes[359:352];
        2029: state_byte <= hashes[351:344];
        2030: state_byte <= hashes[343:336];
        2031: state_byte <= hashes[335:328];
        2032: state_byte <= hashes[327:320];
        2033: state_byte <= hashes[319:312];
        2034: state_byte <= hashes[311:304];
        2035: state_byte <= hashes[303:296];
        2036: state_byte <= hashes[295:288];
        2037: state_byte <= hashes[287:280];
        2038: state_byte <= hashes[279:272];
        2039: state_byte <= hashes[271:264];
        2040: state_byte <= hashes[263:256];
        2041: state_byte <= hashes[255:248];
        2042: state_byte <= hashes[247:240];
        2043: state_byte <= hashes[239:232];
        2044: state_byte <= hashes[231:224];
        2045: state_byte <= hashes[223:216];
        2046: state_byte <= hashes[215:208];
        2047: state_byte <= hashes[207:200];
        2048: state_byte <= hashes[199:192];
        2049: state_byte <= hashes[191:184];
        2050: state_byte <= hashes[183:176];
        2051: state_byte <= hashes[175:168];
        2052: state_byte <= hashes[167:160];
        2053: state_byte <= hashes[159:152];
        2054: state_byte <= hashes[151:144];
        2055: state_byte <= hashes[143:136];
        2056: state_byte <= hashes[135:128];
        2057: state_byte <= hashes[127:120];
        2058: state_byte <= hashes[119:112];
        2059: state_byte <= hashes[111:104];
        2060: state_byte <= hashes[103:96];
        2061: state_byte <= hashes[95:88];
        2062: state_byte <= hashes[87:80];
        2063: state_byte <= hashes[79:72];
        2064: state_byte <= hashes[71:64];
        2065: state_byte <= hashes[63:56];
        2066: state_byte <= hashes[55:48];
        2067: state_byte <= hashes[47:40];
        2068: state_byte <= hashes[39:32];
        2069: state_byte <= hashes[31:24];
        2070: state_byte <= hashes[23:16];
        2071: state_byte <= hashes[15:8];
        2072: state_byte <= hashes[7:0];

        // current hash
        2073: state_byte <= current_hash[127:120];
        2074: state_byte <= current_hash[119:112];
        2075: state_byte <= current_hash[111:104];
        2076: state_byte <= current_hash[103:96];
        2077: state_byte <= current_hash[95:88];
        2078: state_byte <= current_hash[87:80];
        2079: state_byte <= current_hash[79:72];
        2080: state_byte <= current_hash[71:64];
        2081: state_byte <= current_hash[63:56];
        2082: state_byte <= current_hash[55:48];
        2083: state_byte <= current_hash[47:40];
        2084: state_byte <= current_hash[39:32];
        2085: state_byte <= current_hash[31:24];
        2086: state_byte <= current_hash[23:16];
        2087: state_byte <= current_hash[15:8];
        2088: state_byte <= current_hash[7:0];

        // footer
        2089: state_byte <= 8'hA2;
        2090: state_byte <= 8'h5E;
        2091: state_byte <= 8'hFA;
        2092: state_byte <= 8'hCE;

    endcase

    if (byte_index == 2092)
        byte_index <= 0;
    else
        byte_index <= byte_index + 1;
end

endmodule
